VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO systolic_sorter
  CLASS BLOCK ;
  FOREIGN systolic_sorter ;
  ORIGIN 0.000 0.000 ;
  SIZE 1751.000 BY 1751.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 1738.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 1738.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 1738.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 10.640 486.740 1738.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.740 10.640 640.340 1738.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 792.340 10.640 793.940 1738.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 945.940 10.640 947.540 1738.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 1099.540 10.640 1101.140 1738.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 1253.140 10.640 1254.740 1738.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 1406.740 10.640 1408.340 1738.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 1560.340 10.640 1561.940 1738.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 1713.940 10.640 1715.540 1738.320 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 1745.480 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 1745.480 184.810 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 336.390 1745.480 337.990 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 489.570 1745.480 491.170 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 642.750 1745.480 644.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 795.930 1745.480 797.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 949.110 1745.480 950.710 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1102.290 1745.480 1103.890 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1255.470 1745.480 1257.070 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1408.650 1745.480 1410.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1561.830 1745.480 1563.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1715.010 1745.480 1716.610 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1738.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1738.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1738.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1738.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1738.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1738.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1738.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1738.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1738.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1738.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 1738.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 1738.320 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 1745.480 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 1745.480 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 333.090 1745.480 334.690 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 486.270 1745.480 487.870 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 639.450 1745.480 641.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 792.630 1745.480 794.230 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 945.810 1745.480 947.410 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1098.990 1745.480 1100.590 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1252.170 1745.480 1253.770 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1405.350 1745.480 1406.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1558.530 1745.480 1560.130 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1711.710 1745.480 1713.310 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1067.640 4.000 1068.240 ;
    END
  END clk
  PIN in_data_flat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 741.240 1751.000 741.840 ;
    END
  END in_data_flat[0]
  PIN in_data_flat[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1120.650 0.000 1120.930 4.000 ;
    END
  END in_data_flat[100]
  PIN in_data_flat[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1101.330 0.000 1101.610 4.000 ;
    END
  END in_data_flat[101]
  PIN in_data_flat[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1059.470 0.000 1059.750 4.000 ;
    END
  END in_data_flat[102]
  PIN in_data_flat[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1056.250 0.000 1056.530 4.000 ;
    END
  END in_data_flat[103]
  PIN in_data_flat[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 897.640 1751.000 898.240 ;
    END
  END in_data_flat[104]
  PIN in_data_flat[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 928.240 1751.000 928.840 ;
    END
  END in_data_flat[105]
  PIN in_data_flat[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1183.240 1751.000 1183.840 ;
    END
  END in_data_flat[106]
  PIN in_data_flat[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 962.240 1751.000 962.840 ;
    END
  END in_data_flat[107]
  PIN in_data_flat[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1166.240 1751.000 1166.840 ;
    END
  END in_data_flat[108]
  PIN in_data_flat[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1142.440 1751.000 1143.040 ;
    END
  END in_data_flat[109]
  PIN in_data_flat[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 958.840 1751.000 959.440 ;
    END
  END in_data_flat[10]
  PIN in_data_flat[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1159.440 1751.000 1160.040 ;
    END
  END in_data_flat[110]
  PIN in_data_flat[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1084.640 1751.000 1085.240 ;
    END
  END in_data_flat[111]
  PIN in_data_flat[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1009.840 4.000 1010.440 ;
    END
  END in_data_flat[112]
  PIN in_data_flat[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 935.040 4.000 935.640 ;
    END
  END in_data_flat[113]
  PIN in_data_flat[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.240 4.000 758.840 ;
    END
  END in_data_flat[114]
  PIN in_data_flat[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 547.440 4.000 548.040 ;
    END
  END in_data_flat[115]
  PIN in_data_flat[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.040 4.000 561.640 ;
    END
  END in_data_flat[116]
  PIN in_data_flat[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.240 4.000 588.840 ;
    END
  END in_data_flat[117]
  PIN in_data_flat[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END in_data_flat[118]
  PIN in_data_flat[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.840 4.000 721.440 ;
    END
  END in_data_flat[119]
  PIN in_data_flat[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 999.640 1751.000 1000.240 ;
    END
  END in_data_flat[11]
  PIN in_data_flat[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 721.370 1747.000 721.650 1751.000 ;
    END
  END in_data_flat[120]
  PIN in_data_flat[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.040 4.000 884.640 ;
    END
  END in_data_flat[121]
  PIN in_data_flat[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 734.250 1747.000 734.530 1751.000 ;
    END
  END in_data_flat[122]
  PIN in_data_flat[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 737.470 1747.000 737.750 1751.000 ;
    END
  END in_data_flat[123]
  PIN in_data_flat[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 718.150 1747.000 718.430 1751.000 ;
    END
  END in_data_flat[124]
  PIN in_data_flat[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 743.910 1747.000 744.190 1751.000 ;
    END
  END in_data_flat[125]
  PIN in_data_flat[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 747.130 1747.000 747.410 1751.000 ;
    END
  END in_data_flat[126]
  PIN in_data_flat[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 753.570 1747.000 753.850 1751.000 ;
    END
  END in_data_flat[127]
  PIN in_data_flat[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 870.440 1751.000 871.040 ;
    END
  END in_data_flat[128]
  PIN in_data_flat[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 991.850 0.000 992.130 4.000 ;
    END
  END in_data_flat[129]
  PIN in_data_flat[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1040.440 1751.000 1041.040 ;
    END
  END in_data_flat[12]
  PIN in_data_flat[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1014.390 0.000 1014.670 4.000 ;
    END
  END in_data_flat[130]
  PIN in_data_flat[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1027.270 0.000 1027.550 4.000 ;
    END
  END in_data_flat[131]
  PIN in_data_flat[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1078.790 0.000 1079.070 4.000 ;
    END
  END in_data_flat[132]
  PIN in_data_flat[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1007.950 0.000 1008.230 4.000 ;
    END
  END in_data_flat[133]
  PIN in_data_flat[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1017.610 0.000 1017.890 4.000 ;
    END
  END in_data_flat[134]
  PIN in_data_flat[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1020.830 0.000 1021.110 4.000 ;
    END
  END in_data_flat[135]
  PIN in_data_flat[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 890.840 1751.000 891.440 ;
    END
  END in_data_flat[136]
  PIN in_data_flat[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 914.640 1751.000 915.240 ;
    END
  END in_data_flat[137]
  PIN in_data_flat[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1013.240 1751.000 1013.840 ;
    END
  END in_data_flat[138]
  PIN in_data_flat[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 969.040 1751.000 969.640 ;
    END
  END in_data_flat[139]
  PIN in_data_flat[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1135.640 1751.000 1136.240 ;
    END
  END in_data_flat[13]
  PIN in_data_flat[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1118.640 1751.000 1119.240 ;
    END
  END in_data_flat[140]
  PIN in_data_flat[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 995.070 1747.000 995.350 1751.000 ;
    END
  END in_data_flat[141]
  PIN in_data_flat[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1122.040 1751.000 1122.640 ;
    END
  END in_data_flat[142]
  PIN in_data_flat[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1023.440 1751.000 1024.040 ;
    END
  END in_data_flat[143]
  PIN in_data_flat[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 853.440 4.000 854.040 ;
    END
  END in_data_flat[144]
  PIN in_data_flat[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 989.440 4.000 990.040 ;
    END
  END in_data_flat[145]
  PIN in_data_flat[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 761.640 4.000 762.240 ;
    END
  END in_data_flat[146]
  PIN in_data_flat[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.840 4.000 738.440 ;
    END
  END in_data_flat[147]
  PIN in_data_flat[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 4.000 673.840 ;
    END
  END in_data_flat[148]
  PIN in_data_flat[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END in_data_flat[149]
  PIN in_data_flat[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1091.440 1751.000 1092.040 ;
    END
  END in_data_flat[14]
  PIN in_data_flat[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END in_data_flat[150]
  PIN in_data_flat[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.840 4.000 687.440 ;
    END
  END in_data_flat[151]
  PIN in_data_flat[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 901.040 4.000 901.640 ;
    END
  END in_data_flat[152]
  PIN in_data_flat[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 873.840 4.000 874.440 ;
    END
  END in_data_flat[153]
  PIN in_data_flat[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 986.040 4.000 986.640 ;
    END
  END in_data_flat[154]
  PIN in_data_flat[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 695.610 1747.000 695.890 1751.000 ;
    END
  END in_data_flat[155]
  PIN in_data_flat[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 698.830 1747.000 699.110 1751.000 ;
    END
  END in_data_flat[156]
  PIN in_data_flat[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 702.050 1747.000 702.330 1751.000 ;
    END
  END in_data_flat[157]
  PIN in_data_flat[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 692.390 1747.000 692.670 1751.000 ;
    END
  END in_data_flat[158]
  PIN in_data_flat[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 705.270 1747.000 705.550 1751.000 ;
    END
  END in_data_flat[159]
  PIN in_data_flat[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1020.040 1751.000 1020.640 ;
    END
  END in_data_flat[15]
  PIN in_data_flat[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 969.310 0.000 969.590 4.000 ;
    END
  END in_data_flat[160]
  PIN in_data_flat[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 959.650 0.000 959.930 4.000 ;
    END
  END in_data_flat[161]
  PIN in_data_flat[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 972.530 0.000 972.810 4.000 ;
    END
  END in_data_flat[162]
  PIN in_data_flat[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 962.870 0.000 963.150 4.000 ;
    END
  END in_data_flat[163]
  PIN in_data_flat[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 982.190 0.000 982.470 4.000 ;
    END
  END in_data_flat[164]
  PIN in_data_flat[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 956.430 0.000 956.710 4.000 ;
    END
  END in_data_flat[165]
  PIN in_data_flat[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 978.970 0.000 979.250 4.000 ;
    END
  END in_data_flat[166]
  PIN in_data_flat[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 975.750 0.000 976.030 4.000 ;
    END
  END in_data_flat[167]
  PIN in_data_flat[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 966.090 0.000 966.370 4.000 ;
    END
  END in_data_flat[168]
  PIN in_data_flat[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 765.040 1751.000 765.640 ;
    END
  END in_data_flat[169]
  PIN in_data_flat[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 760.010 0.000 760.290 4.000 ;
    END
  END in_data_flat[16]
  PIN in_data_flat[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 989.440 1751.000 990.040 ;
    END
  END in_data_flat[170]
  PIN in_data_flat[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 955.440 1751.000 956.040 ;
    END
  END in_data_flat[171]
  PIN in_data_flat[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1064.240 1751.000 1064.840 ;
    END
  END in_data_flat[172]
  PIN in_data_flat[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 969.310 1747.000 969.590 1751.000 ;
    END
  END in_data_flat[173]
  PIN in_data_flat[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 966.090 1747.000 966.370 1751.000 ;
    END
  END in_data_flat[174]
  PIN in_data_flat[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1016.640 1751.000 1017.240 ;
    END
  END in_data_flat[175]
  PIN in_data_flat[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.240 4.000 843.840 ;
    END
  END in_data_flat[176]
  PIN in_data_flat[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 833.040 4.000 833.640 ;
    END
  END in_data_flat[177]
  PIN in_data_flat[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 768.440 4.000 769.040 ;
    END
  END in_data_flat[178]
  PIN in_data_flat[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.040 4.000 646.640 ;
    END
  END in_data_flat[179]
  PIN in_data_flat[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 850.170 0.000 850.450 4.000 ;
    END
  END in_data_flat[17]
  PIN in_data_flat[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END in_data_flat[180]
  PIN in_data_flat[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END in_data_flat[181]
  PIN in_data_flat[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.840 4.000 670.440 ;
    END
  END in_data_flat[182]
  PIN in_data_flat[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.040 4.000 714.640 ;
    END
  END in_data_flat[183]
  PIN in_data_flat[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 894.240 4.000 894.840 ;
    END
  END in_data_flat[184]
  PIN in_data_flat[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 870.440 4.000 871.040 ;
    END
  END in_data_flat[185]
  PIN in_data_flat[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 941.840 4.000 942.440 ;
    END
  END in_data_flat[186]
  PIN in_data_flat[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 982.640 4.000 983.240 ;
    END
  END in_data_flat[187]
  PIN in_data_flat[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 656.970 1747.000 657.250 1751.000 ;
    END
  END in_data_flat[188]
  PIN in_data_flat[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 660.190 1747.000 660.470 1751.000 ;
    END
  END in_data_flat[189]
  PIN in_data_flat[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 859.830 0.000 860.110 4.000 ;
    END
  END in_data_flat[18]
  PIN in_data_flat[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 666.630 1747.000 666.910 1751.000 ;
    END
  END in_data_flat[190]
  PIN in_data_flat[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 673.070 1747.000 673.350 1751.000 ;
    END
  END in_data_flat[191]
  PIN in_data_flat[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 930.670 0.000 930.950 4.000 ;
    END
  END in_data_flat[192]
  PIN in_data_flat[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 898.470 0.000 898.750 4.000 ;
    END
  END in_data_flat[193]
  PIN in_data_flat[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 924.230 0.000 924.510 4.000 ;
    END
  END in_data_flat[194]
  PIN in_data_flat[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 914.570 0.000 914.850 4.000 ;
    END
  END in_data_flat[195]
  PIN in_data_flat[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 785.770 0.000 786.050 4.000 ;
    END
  END in_data_flat[196]
  PIN in_data_flat[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 917.790 0.000 918.070 4.000 ;
    END
  END in_data_flat[197]
  PIN in_data_flat[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 937.110 0.000 937.390 4.000 ;
    END
  END in_data_flat[198]
  PIN in_data_flat[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 940.330 0.000 940.610 4.000 ;
    END
  END in_data_flat[199]
  PIN in_data_flat[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 853.390 0.000 853.670 4.000 ;
    END
  END in_data_flat[19]
  PIN in_data_flat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 843.240 1751.000 843.840 ;
    END
  END in_data_flat[1]
  PIN in_data_flat[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 921.010 0.000 921.290 4.000 ;
    END
  END in_data_flat[200]
  PIN in_data_flat[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 927.450 0.000 927.730 4.000 ;
    END
  END in_data_flat[201]
  PIN in_data_flat[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 975.840 1751.000 976.440 ;
    END
  END in_data_flat[202]
  PIN in_data_flat[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 952.040 1751.000 952.640 ;
    END
  END in_data_flat[203]
  PIN in_data_flat[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 946.770 1747.000 947.050 1751.000 ;
    END
  END in_data_flat[204]
  PIN in_data_flat[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 921.010 1747.000 921.290 1751.000 ;
    END
  END in_data_flat[205]
  PIN in_data_flat[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 914.570 1747.000 914.850 1751.000 ;
    END
  END in_data_flat[206]
  PIN in_data_flat[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1003.040 1751.000 1003.640 ;
    END
  END in_data_flat[207]
  PIN in_data_flat[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 931.640 4.000 932.240 ;
    END
  END in_data_flat[208]
  PIN in_data_flat[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1003.040 4.000 1003.640 ;
    END
  END in_data_flat[209]
  PIN in_data_flat[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 843.730 0.000 844.010 4.000 ;
    END
  END in_data_flat[20]
  PIN in_data_flat[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.040 4.000 765.640 ;
    END
  END in_data_flat[210]
  PIN in_data_flat[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END in_data_flat[211]
  PIN in_data_flat[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END in_data_flat[212]
  PIN in_data_flat[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 608.640 4.000 609.240 ;
    END
  END in_data_flat[213]
  PIN in_data_flat[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.040 4.000 663.640 ;
    END
  END in_data_flat[214]
  PIN in_data_flat[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.240 4.000 571.840 ;
    END
  END in_data_flat[215]
  PIN in_data_flat[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 887.440 4.000 888.040 ;
    END
  END in_data_flat[216]
  PIN in_data_flat[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 860.240 4.000 860.840 ;
    END
  END in_data_flat[217]
  PIN in_data_flat[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 962.240 4.000 962.840 ;
    END
  END in_data_flat[218]
  PIN in_data_flat[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 969.040 4.000 969.640 ;
    END
  END in_data_flat[219]
  PIN in_data_flat[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 846.950 0.000 847.230 4.000 ;
    END
  END in_data_flat[21]
  PIN in_data_flat[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 647.310 1747.000 647.590 1751.000 ;
    END
  END in_data_flat[220]
  PIN in_data_flat[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 634.430 1747.000 634.710 1751.000 ;
    END
  END in_data_flat[221]
  PIN in_data_flat[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1020.040 4.000 1020.640 ;
    END
  END in_data_flat[222]
  PIN in_data_flat[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 996.240 4.000 996.840 ;
    END
  END in_data_flat[223]
  PIN in_data_flat[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 888.810 0.000 889.090 4.000 ;
    END
  END in_data_flat[224]
  PIN in_data_flat[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 866.270 0.000 866.550 4.000 ;
    END
  END in_data_flat[225]
  PIN in_data_flat[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 840.510 0.000 840.790 4.000 ;
    END
  END in_data_flat[226]
  PIN in_data_flat[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 872.710 0.000 872.990 4.000 ;
    END
  END in_data_flat[227]
  PIN in_data_flat[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 782.550 0.000 782.830 4.000 ;
    END
  END in_data_flat[228]
  PIN in_data_flat[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 875.930 0.000 876.210 4.000 ;
    END
  END in_data_flat[229]
  PIN in_data_flat[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 856.610 0.000 856.890 4.000 ;
    END
  END in_data_flat[22]
  PIN in_data_flat[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 904.910 0.000 905.190 4.000 ;
    END
  END in_data_flat[230]
  PIN in_data_flat[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 901.690 0.000 901.970 4.000 ;
    END
  END in_data_flat[231]
  PIN in_data_flat[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 788.990 0.000 789.270 4.000 ;
    END
  END in_data_flat[232]
  PIN in_data_flat[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 924.230 1747.000 924.510 1751.000 ;
    END
  END in_data_flat[233]
  PIN in_data_flat[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 888.810 1747.000 889.090 1751.000 ;
    END
  END in_data_flat[234]
  PIN in_data_flat[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 927.450 1747.000 927.730 1751.000 ;
    END
  END in_data_flat[235]
  PIN in_data_flat[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 875.930 1747.000 876.210 1751.000 ;
    END
  END in_data_flat[236]
  PIN in_data_flat[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 892.030 1747.000 892.310 1751.000 ;
    END
  END in_data_flat[237]
  PIN in_data_flat[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 885.590 1747.000 885.870 1751.000 ;
    END
  END in_data_flat[238]
  PIN in_data_flat[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 882.370 1747.000 882.650 1751.000 ;
    END
  END in_data_flat[239]
  PIN in_data_flat[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 863.050 0.000 863.330 4.000 ;
    END
  END in_data_flat[23]
  PIN in_data_flat[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.840 4.000 840.440 ;
    END
  END in_data_flat[240]
  PIN in_data_flat[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 809.240 4.000 809.840 ;
    END
  END in_data_flat[241]
  PIN in_data_flat[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.040 4.000 782.640 ;
    END
  END in_data_flat[242]
  PIN in_data_flat[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 754.840 4.000 755.440 ;
    END
  END in_data_flat[243]
  PIN in_data_flat[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 649.440 4.000 650.040 ;
    END
  END in_data_flat[244]
  PIN in_data_flat[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.040 4.000 595.640 ;
    END
  END in_data_flat[245]
  PIN in_data_flat[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END in_data_flat[246]
  PIN in_data_flat[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.040 4.000 731.640 ;
    END
  END in_data_flat[247]
  PIN in_data_flat[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 890.840 4.000 891.440 ;
    END
  END in_data_flat[248]
  PIN in_data_flat[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 863.640 4.000 864.240 ;
    END
  END in_data_flat[249]
  PIN in_data_flat[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 956.430 1747.000 956.710 1751.000 ;
    END
  END in_data_flat[24]
  PIN in_data_flat[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 914.640 4.000 915.240 ;
    END
  END in_data_flat[250]
  PIN in_data_flat[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 979.240 4.000 979.840 ;
    END
  END in_data_flat[251]
  PIN in_data_flat[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 621.550 1747.000 621.830 1751.000 ;
    END
  END in_data_flat[252]
  PIN in_data_flat[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 618.330 1747.000 618.610 1751.000 ;
    END
  END in_data_flat[253]
  PIN in_data_flat[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 595.790 1747.000 596.070 1751.000 ;
    END
  END in_data_flat[254]
  PIN in_data_flat[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 992.840 4.000 993.440 ;
    END
  END in_data_flat[255]
  PIN in_data_flat[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 859.830 1747.000 860.110 1751.000 ;
    END
  END in_data_flat[25]
  PIN in_data_flat[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 872.710 1747.000 872.990 1751.000 ;
    END
  END in_data_flat[26]
  PIN in_data_flat[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 953.210 1747.000 953.490 1751.000 ;
    END
  END in_data_flat[27]
  PIN in_data_flat[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 940.330 1747.000 940.610 1751.000 ;
    END
  END in_data_flat[28]
  PIN in_data_flat[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 856.610 1747.000 856.890 1751.000 ;
    END
  END in_data_flat[29]
  PIN in_data_flat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 805.840 1751.000 806.440 ;
    END
  END in_data_flat[2]
  PIN in_data_flat[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 853.390 1747.000 853.670 1751.000 ;
    END
  END in_data_flat[30]
  PIN in_data_flat[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 840.510 1747.000 840.790 1751.000 ;
    END
  END in_data_flat[31]
  PIN in_data_flat[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 877.240 1751.000 877.840 ;
    END
  END in_data_flat[32]
  PIN in_data_flat[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 850.040 1751.000 850.640 ;
    END
  END in_data_flat[33]
  PIN in_data_flat[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 809.240 1751.000 809.840 ;
    END
  END in_data_flat[34]
  PIN in_data_flat[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 782.040 1751.000 782.640 ;
    END
  END in_data_flat[35]
  PIN in_data_flat[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1133.530 0.000 1133.810 4.000 ;
    END
  END in_data_flat[36]
  PIN in_data_flat[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1130.310 0.000 1130.590 4.000 ;
    END
  END in_data_flat[37]
  PIN in_data_flat[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 720.840 1751.000 721.440 ;
    END
  END in_data_flat[38]
  PIN in_data_flat[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 744.640 1751.000 745.240 ;
    END
  END in_data_flat[39]
  PIN in_data_flat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 795.640 1751.000 796.240 ;
    END
  END in_data_flat[3]
  PIN in_data_flat[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 901.040 1751.000 901.640 ;
    END
  END in_data_flat[40]
  PIN in_data_flat[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 918.040 1751.000 918.640 ;
    END
  END in_data_flat[41]
  PIN in_data_flat[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 965.640 1751.000 966.240 ;
    END
  END in_data_flat[42]
  PIN in_data_flat[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 992.840 1751.000 993.440 ;
    END
  END in_data_flat[43]
  PIN in_data_flat[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1149.240 1751.000 1149.840 ;
    END
  END in_data_flat[44]
  PIN in_data_flat[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1105.040 1751.000 1105.640 ;
    END
  END in_data_flat[45]
  PIN in_data_flat[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1179.840 1751.000 1180.440 ;
    END
  END in_data_flat[46]
  PIN in_data_flat[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1026.840 1751.000 1027.440 ;
    END
  END in_data_flat[47]
  PIN in_data_flat[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 850.040 4.000 850.640 ;
    END
  END in_data_flat[48]
  PIN in_data_flat[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 829.640 4.000 830.240 ;
    END
  END in_data_flat[49]
  PIN in_data_flat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1152.850 0.000 1153.130 4.000 ;
    END
  END in_data_flat[4]
  PIN in_data_flat[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 775.240 4.000 775.840 ;
    END
  END in_data_flat[50]
  PIN in_data_flat[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 748.040 4.000 748.640 ;
    END
  END in_data_flat[51]
  PIN in_data_flat[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 805.090 0.000 805.370 4.000 ;
    END
  END in_data_flat[52]
  PIN in_data_flat[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 814.750 0.000 815.030 4.000 ;
    END
  END in_data_flat[53]
  PIN in_data_flat[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 827.630 0.000 827.910 4.000 ;
    END
  END in_data_flat[54]
  PIN in_data_flat[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 727.640 4.000 728.240 ;
    END
  END in_data_flat[55]
  PIN in_data_flat[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 837.290 1747.000 837.570 1751.000 ;
    END
  END in_data_flat[56]
  PIN in_data_flat[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 817.970 1747.000 818.250 1751.000 ;
    END
  END in_data_flat[57]
  PIN in_data_flat[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 821.190 1747.000 821.470 1751.000 ;
    END
  END in_data_flat[58]
  PIN in_data_flat[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 843.730 1747.000 844.010 1751.000 ;
    END
  END in_data_flat[59]
  PIN in_data_flat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1127.090 0.000 1127.370 4.000 ;
    END
  END in_data_flat[5]
  PIN in_data_flat[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 834.070 1747.000 834.350 1751.000 ;
    END
  END in_data_flat[60]
  PIN in_data_flat[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 830.850 1747.000 831.130 1751.000 ;
    END
  END in_data_flat[61]
  PIN in_data_flat[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 827.630 1747.000 827.910 1751.000 ;
    END
  END in_data_flat[62]
  PIN in_data_flat[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 824.410 1747.000 824.690 1751.000 ;
    END
  END in_data_flat[63]
  PIN in_data_flat[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 867.040 1751.000 867.640 ;
    END
  END in_data_flat[64]
  PIN in_data_flat[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 846.640 1751.000 847.240 ;
    END
  END in_data_flat[65]
  PIN in_data_flat[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 819.440 1751.000 820.040 ;
    END
  END in_data_flat[66]
  PIN in_data_flat[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 792.240 1751.000 792.840 ;
    END
  END in_data_flat[67]
  PIN in_data_flat[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1091.670 0.000 1091.950 4.000 ;
    END
  END in_data_flat[68]
  PIN in_data_flat[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1098.110 0.000 1098.390 4.000 ;
    END
  END in_data_flat[69]
  PIN in_data_flat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 737.840 1751.000 738.440 ;
    END
  END in_data_flat[6]
  PIN in_data_flat[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1088.450 0.000 1088.730 4.000 ;
    END
  END in_data_flat[70]
  PIN in_data_flat[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1094.890 0.000 1095.170 4.000 ;
    END
  END in_data_flat[71]
  PIN in_data_flat[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 880.640 1751.000 881.240 ;
    END
  END in_data_flat[72]
  PIN in_data_flat[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 924.840 1751.000 925.440 ;
    END
  END in_data_flat[73]
  PIN in_data_flat[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 979.240 1751.000 979.840 ;
    END
  END in_data_flat[74]
  PIN in_data_flat[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1043.840 1751.000 1044.440 ;
    END
  END in_data_flat[75]
  PIN in_data_flat[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1125.440 1751.000 1126.040 ;
    END
  END in_data_flat[76]
  PIN in_data_flat[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1128.840 1751.000 1129.440 ;
    END
  END in_data_flat[77]
  PIN in_data_flat[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1169.640 1751.000 1170.240 ;
    END
  END in_data_flat[78]
  PIN in_data_flat[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1009.840 1751.000 1010.440 ;
    END
  END in_data_flat[79]
  PIN in_data_flat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 771.840 1751.000 772.440 ;
    END
  END in_data_flat[7]
  PIN in_data_flat[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 897.640 4.000 898.240 ;
    END
  END in_data_flat[80]
  PIN in_data_flat[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 819.440 4.000 820.040 ;
    END
  END in_data_flat[81]
  PIN in_data_flat[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 771.840 4.000 772.440 ;
    END
  END in_data_flat[82]
  PIN in_data_flat[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.040 4.000 697.640 ;
    END
  END in_data_flat[83]
  PIN in_data_flat[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.240 4.000 622.840 ;
    END
  END in_data_flat[84]
  PIN in_data_flat[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 779.330 0.000 779.610 4.000 ;
    END
  END in_data_flat[85]
  PIN in_data_flat[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 776.110 0.000 776.390 4.000 ;
    END
  END in_data_flat[86]
  PIN in_data_flat[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.840 4.000 568.440 ;
    END
  END in_data_flat[87]
  PIN in_data_flat[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 788.990 1747.000 789.270 1751.000 ;
    END
  END in_data_flat[88]
  PIN in_data_flat[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 785.770 1747.000 786.050 1751.000 ;
    END
  END in_data_flat[89]
  PIN in_data_flat[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 904.440 1751.000 905.040 ;
    END
  END in_data_flat[8]
  PIN in_data_flat[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 769.670 1747.000 769.950 1751.000 ;
    END
  END in_data_flat[90]
  PIN in_data_flat[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 772.890 1747.000 773.170 1751.000 ;
    END
  END in_data_flat[91]
  PIN in_data_flat[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 798.650 1747.000 798.930 1751.000 ;
    END
  END in_data_flat[92]
  PIN in_data_flat[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 782.550 1747.000 782.830 1751.000 ;
    END
  END in_data_flat[93]
  PIN in_data_flat[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 779.330 1747.000 779.610 1751.000 ;
    END
  END in_data_flat[94]
  PIN in_data_flat[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 776.110 1747.000 776.390 1751.000 ;
    END
  END in_data_flat[95]
  PIN in_data_flat[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 826.240 1751.000 826.840 ;
    END
  END in_data_flat[96]
  PIN in_data_flat[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 853.440 1751.000 854.040 ;
    END
  END in_data_flat[97]
  PIN in_data_flat[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1043.370 0.000 1043.650 4.000 ;
    END
  END in_data_flat[98]
  PIN in_data_flat[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1075.570 0.000 1075.850 4.000 ;
    END
  END in_data_flat[99]
  PIN in_data_flat[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 931.640 1751.000 932.240 ;
    END
  END in_data_flat[9]
  PIN load
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1064.240 4.000 1064.840 ;
    END
  END load
  PIN out_data_flat[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 860.240 1751.000 860.840 ;
    END
  END out_data_flat[0]
  PIN out_data_flat[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1082.010 0.000 1082.290 4.000 ;
    END
  END out_data_flat[100]
  PIN out_data_flat[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1104.550 0.000 1104.830 4.000 ;
    END
  END out_data_flat[101]
  PIN out_data_flat[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1072.350 0.000 1072.630 4.000 ;
    END
  END out_data_flat[102]
  PIN out_data_flat[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1085.230 0.000 1085.510 4.000 ;
    END
  END out_data_flat[103]
  PIN out_data_flat[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 884.040 1751.000 884.640 ;
    END
  END out_data_flat[104]
  PIN out_data_flat[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 921.440 1751.000 922.040 ;
    END
  END out_data_flat[105]
  PIN out_data_flat[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1057.440 1751.000 1058.040 ;
    END
  END out_data_flat[106]
  PIN out_data_flat[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 972.440 1751.000 973.040 ;
    END
  END out_data_flat[107]
  PIN out_data_flat[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1077.840 1751.000 1078.440 ;
    END
  END out_data_flat[108]
  PIN out_data_flat[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1132.240 1751.000 1132.840 ;
    END
  END out_data_flat[109]
  PIN out_data_flat[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 941.840 1751.000 942.440 ;
    END
  END out_data_flat[10]
  PIN out_data_flat[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1145.840 1751.000 1146.440 ;
    END
  END out_data_flat[110]
  PIN out_data_flat[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1054.040 1751.000 1054.640 ;
    END
  END out_data_flat[111]
  PIN out_data_flat[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 904.440 4.000 905.040 ;
    END
  END out_data_flat[112]
  PIN out_data_flat[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 816.040 4.000 816.640 ;
    END
  END out_data_flat[113]
  PIN out_data_flat[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 778.640 4.000 779.240 ;
    END
  END out_data_flat[114]
  PIN out_data_flat[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 744.640 4.000 745.240 ;
    END
  END out_data_flat[115]
  PIN out_data_flat[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 676.640 4.000 677.240 ;
    END
  END out_data_flat[116]
  PIN out_data_flat[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.040 4.000 629.640 ;
    END
  END out_data_flat[117]
  PIN out_data_flat[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.840 4.000 636.440 ;
    END
  END out_data_flat[118]
  PIN out_data_flat[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.240 4.000 690.840 ;
    END
  END out_data_flat[119]
  PIN out_data_flat[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 986.040 1751.000 986.640 ;
    END
  END out_data_flat[11]
  PIN out_data_flat[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 714.930 1747.000 715.210 1751.000 ;
    END
  END out_data_flat[120]
  PIN out_data_flat[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 724.590 1747.000 724.870 1751.000 ;
    END
  END out_data_flat[121]
  PIN out_data_flat[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 682.730 1747.000 683.010 1751.000 ;
    END
  END out_data_flat[122]
  PIN out_data_flat[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 711.710 1747.000 711.990 1751.000 ;
    END
  END out_data_flat[123]
  PIN out_data_flat[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 685.950 1747.000 686.230 1751.000 ;
    END
  END out_data_flat[124]
  PIN out_data_flat[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 708.490 1747.000 708.770 1751.000 ;
    END
  END out_data_flat[125]
  PIN out_data_flat[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 727.810 1747.000 728.090 1751.000 ;
    END
  END out_data_flat[126]
  PIN out_data_flat[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 689.170 1747.000 689.450 1751.000 ;
    END
  END out_data_flat[127]
  PIN out_data_flat[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1062.690 0.000 1062.970 4.000 ;
    END
  END out_data_flat[128]
  PIN out_data_flat[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1053.030 0.000 1053.310 4.000 ;
    END
  END out_data_flat[129]
  PIN out_data_flat[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1060.840 1751.000 1061.440 ;
    END
  END out_data_flat[12]
  PIN out_data_flat[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1036.930 0.000 1037.210 4.000 ;
    END
  END out_data_flat[130]
  PIN out_data_flat[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1046.590 0.000 1046.870 4.000 ;
    END
  END out_data_flat[131]
  PIN out_data_flat[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1040.150 0.000 1040.430 4.000 ;
    END
  END out_data_flat[132]
  PIN out_data_flat[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1033.710 0.000 1033.990 4.000 ;
    END
  END out_data_flat[133]
  PIN out_data_flat[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1030.490 0.000 1030.770 4.000 ;
    END
  END out_data_flat[134]
  PIN out_data_flat[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1049.810 0.000 1050.090 4.000 ;
    END
  END out_data_flat[135]
  PIN out_data_flat[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 887.440 1751.000 888.040 ;
    END
  END out_data_flat[136]
  PIN out_data_flat[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 911.240 1751.000 911.840 ;
    END
  END out_data_flat[137]
  PIN out_data_flat[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1067.640 1751.000 1068.240 ;
    END
  END out_data_flat[138]
  PIN out_data_flat[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 948.640 1751.000 949.240 ;
    END
  END out_data_flat[139]
  PIN out_data_flat[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1094.840 1751.000 1095.440 ;
    END
  END out_data_flat[13]
  PIN out_data_flat[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1173.040 1751.000 1173.640 ;
    END
  END out_data_flat[140]
  PIN out_data_flat[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1115.240 1751.000 1115.840 ;
    END
  END out_data_flat[141]
  PIN out_data_flat[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1152.640 1751.000 1153.240 ;
    END
  END out_data_flat[142]
  PIN out_data_flat[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1047.240 1751.000 1047.840 ;
    END
  END out_data_flat[143]
  PIN out_data_flat[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 846.640 4.000 847.240 ;
    END
  END out_data_flat[144]
  PIN out_data_flat[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1006.440 4.000 1007.040 ;
    END
  END out_data_flat[145]
  PIN out_data_flat[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 802.440 4.000 803.040 ;
    END
  END out_data_flat[146]
  PIN out_data_flat[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 734.440 4.000 735.040 ;
    END
  END out_data_flat[147]
  PIN out_data_flat[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END out_data_flat[148]
  PIN out_data_flat[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END out_data_flat[149]
  PIN out_data_flat[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1074.440 1751.000 1075.040 ;
    END
  END out_data_flat[14]
  PIN out_data_flat[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.840 4.000 602.440 ;
    END
  END out_data_flat[150]
  PIN out_data_flat[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END out_data_flat[151]
  PIN out_data_flat[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 952.040 4.000 952.640 ;
    END
  END out_data_flat[152]
  PIN out_data_flat[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 958.840 4.000 959.440 ;
    END
  END out_data_flat[153]
  PIN out_data_flat[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 948.640 4.000 949.240 ;
    END
  END out_data_flat[154]
  PIN out_data_flat[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 663.410 1747.000 663.690 1751.000 ;
    END
  END out_data_flat[155]
  PIN out_data_flat[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 676.290 1747.000 676.570 1751.000 ;
    END
  END out_data_flat[156]
  PIN out_data_flat[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 669.850 1747.000 670.130 1751.000 ;
    END
  END out_data_flat[157]
  PIN out_data_flat[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 679.510 1747.000 679.790 1751.000 ;
    END
  END out_data_flat[158]
  PIN out_data_flat[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 653.750 1747.000 654.030 1751.000 ;
    END
  END out_data_flat[159]
  PIN out_data_flat[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1030.240 1751.000 1030.840 ;
    END
  END out_data_flat[15]
  PIN out_data_flat[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 988.630 0.000 988.910 4.000 ;
    END
  END out_data_flat[160]
  PIN out_data_flat[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 998.290 0.000 998.570 4.000 ;
    END
  END out_data_flat[161]
  PIN out_data_flat[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 995.070 0.000 995.350 4.000 ;
    END
  END out_data_flat[162]
  PIN out_data_flat[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1004.730 0.000 1005.010 4.000 ;
    END
  END out_data_flat[163]
  PIN out_data_flat[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1001.510 0.000 1001.790 4.000 ;
    END
  END out_data_flat[164]
  PIN out_data_flat[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 985.410 0.000 985.690 4.000 ;
    END
  END out_data_flat[165]
  PIN out_data_flat[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1024.050 0.000 1024.330 4.000 ;
    END
  END out_data_flat[166]
  PIN out_data_flat[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1011.170 0.000 1011.450 4.000 ;
    END
  END out_data_flat[167]
  PIN out_data_flat[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 856.840 1751.000 857.440 ;
    END
  END out_data_flat[168]
  PIN out_data_flat[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 761.640 1751.000 762.240 ;
    END
  END out_data_flat[169]
  PIN out_data_flat[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 817.970 0.000 818.250 4.000 ;
    END
  END out_data_flat[16]
  PIN out_data_flat[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1006.440 1751.000 1007.040 ;
    END
  END out_data_flat[170]
  PIN out_data_flat[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 938.440 1751.000 939.040 ;
    END
  END out_data_flat[171]
  PIN out_data_flat[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1081.240 1751.000 1081.840 ;
    END
  END out_data_flat[172]
  PIN out_data_flat[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1156.040 1751.000 1156.640 ;
    END
  END out_data_flat[173]
  PIN out_data_flat[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1176.440 1751.000 1177.040 ;
    END
  END out_data_flat[174]
  PIN out_data_flat[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1037.040 1751.000 1037.640 ;
    END
  END out_data_flat[175]
  PIN out_data_flat[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 907.840 4.000 908.440 ;
    END
  END out_data_flat[176]
  PIN out_data_flat[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 999.640 4.000 1000.240 ;
    END
  END out_data_flat[177]
  PIN out_data_flat[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.040 4.000 799.640 ;
    END
  END out_data_flat[178]
  PIN out_data_flat[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END out_data_flat[179]
  PIN out_data_flat[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 824.410 0.000 824.690 4.000 ;
    END
  END out_data_flat[17]
  PIN out_data_flat[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 656.240 4.000 656.840 ;
    END
  END out_data_flat[180]
  PIN out_data_flat[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 615.440 4.000 616.040 ;
    END
  END out_data_flat[181]
  PIN out_data_flat[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END out_data_flat[182]
  PIN out_data_flat[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.240 4.000 707.840 ;
    END
  END out_data_flat[183]
  PIN out_data_flat[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 918.040 4.000 918.640 ;
    END
  END out_data_flat[184]
  PIN out_data_flat[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 880.640 4.000 881.240 ;
    END
  END out_data_flat[185]
  PIN out_data_flat[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 945.240 4.000 945.840 ;
    END
  END out_data_flat[186]
  PIN out_data_flat[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 975.840 4.000 976.440 ;
    END
  END out_data_flat[187]
  PIN out_data_flat[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 650.530 1747.000 650.810 1751.000 ;
    END
  END out_data_flat[188]
  PIN out_data_flat[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 644.090 1747.000 644.370 1751.000 ;
    END
  END out_data_flat[189]
  PIN out_data_flat[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 830.850 0.000 831.130 4.000 ;
    END
  END out_data_flat[18]
  PIN out_data_flat[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 637.650 1747.000 637.930 1751.000 ;
    END
  END out_data_flat[190]
  PIN out_data_flat[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 640.870 1747.000 641.150 1751.000 ;
    END
  END out_data_flat[191]
  PIN out_data_flat[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 895.250 0.000 895.530 4.000 ;
    END
  END out_data_flat[192]
  PIN out_data_flat[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 792.210 0.000 792.490 4.000 ;
    END
  END out_data_flat[193]
  PIN out_data_flat[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 933.890 0.000 934.170 4.000 ;
    END
  END out_data_flat[194]
  PIN out_data_flat[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 943.550 0.000 943.830 4.000 ;
    END
  END out_data_flat[195]
  PIN out_data_flat[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 772.890 0.000 773.170 4.000 ;
    END
  END out_data_flat[196]
  PIN out_data_flat[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 885.590 0.000 885.870 4.000 ;
    END
  END out_data_flat[197]
  PIN out_data_flat[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 946.770 0.000 947.050 4.000 ;
    END
  END out_data_flat[198]
  PIN out_data_flat[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 953.210 0.000 953.490 4.000 ;
    END
  END out_data_flat[199]
  PIN out_data_flat[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 834.070 0.000 834.350 4.000 ;
    END
  END out_data_flat[19]
  PIN out_data_flat[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 839.840 1751.000 840.440 ;
    END
  END out_data_flat[1]
  PIN out_data_flat[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 949.990 0.000 950.270 4.000 ;
    END
  END out_data_flat[200]
  PIN out_data_flat[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 894.240 1751.000 894.840 ;
    END
  END out_data_flat[201]
  PIN out_data_flat[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 935.040 1751.000 935.640 ;
    END
  END out_data_flat[202]
  PIN out_data_flat[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 751.440 1751.000 752.040 ;
    END
  END out_data_flat[203]
  PIN out_data_flat[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 933.890 1747.000 934.170 1751.000 ;
    END
  END out_data_flat[204]
  PIN out_data_flat[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 943.550 1747.000 943.830 1751.000 ;
    END
  END out_data_flat[205]
  PIN out_data_flat[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 930.670 1747.000 930.950 1751.000 ;
    END
  END out_data_flat[206]
  PIN out_data_flat[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1033.640 1751.000 1034.240 ;
    END
  END out_data_flat[207]
  PIN out_data_flat[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 928.240 4.000 928.840 ;
    END
  END out_data_flat[208]
  PIN out_data_flat[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 805.840 4.000 806.440 ;
    END
  END out_data_flat[209]
  PIN out_data_flat[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 811.530 0.000 811.810 4.000 ;
    END
  END out_data_flat[20]
  PIN out_data_flat[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.840 4.000 789.440 ;
    END
  END out_data_flat[210]
  PIN out_data_flat[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 724.240 4.000 724.840 ;
    END
  END out_data_flat[211]
  PIN out_data_flat[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.240 4.000 554.840 ;
    END
  END out_data_flat[212]
  PIN out_data_flat[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.040 4.000 612.640 ;
    END
  END out_data_flat[213]
  PIN out_data_flat[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 683.440 4.000 684.040 ;
    END
  END out_data_flat[214]
  PIN out_data_flat[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END out_data_flat[215]
  PIN out_data_flat[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 911.240 4.000 911.840 ;
    END
  END out_data_flat[216]
  PIN out_data_flat[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 924.840 4.000 925.440 ;
    END
  END out_data_flat[217]
  PIN out_data_flat[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 955.440 4.000 956.040 ;
    END
  END out_data_flat[218]
  PIN out_data_flat[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 972.440 4.000 973.040 ;
    END
  END out_data_flat[219]
  PIN out_data_flat[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 808.310 0.000 808.590 4.000 ;
    END
  END out_data_flat[21]
  PIN out_data_flat[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 631.210 1747.000 631.490 1751.000 ;
    END
  END out_data_flat[220]
  PIN out_data_flat[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 627.990 1747.000 628.270 1751.000 ;
    END
  END out_data_flat[221]
  PIN out_data_flat[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 608.670 1747.000 608.950 1751.000 ;
    END
  END out_data_flat[222]
  PIN out_data_flat[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 611.890 1747.000 612.170 1751.000 ;
    END
  END out_data_flat[223]
  PIN out_data_flat[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 892.030 0.000 892.310 4.000 ;
    END
  END out_data_flat[224]
  PIN out_data_flat[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 879.150 0.000 879.430 4.000 ;
    END
  END out_data_flat[225]
  PIN out_data_flat[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 766.450 0.000 766.730 4.000 ;
    END
  END out_data_flat[226]
  PIN out_data_flat[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 882.370 0.000 882.650 4.000 ;
    END
  END out_data_flat[227]
  PIN out_data_flat[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 769.670 0.000 769.950 4.000 ;
    END
  END out_data_flat[228]
  PIN out_data_flat[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 869.490 0.000 869.770 4.000 ;
    END
  END out_data_flat[229]
  PIN out_data_flat[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 821.190 0.000 821.470 4.000 ;
    END
  END out_data_flat[22]
  PIN out_data_flat[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 908.130 0.000 908.410 4.000 ;
    END
  END out_data_flat[230]
  PIN out_data_flat[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 911.350 0.000 911.630 4.000 ;
    END
  END out_data_flat[231]
  PIN out_data_flat[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 763.230 0.000 763.510 4.000 ;
    END
  END out_data_flat[232]
  PIN out_data_flat[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 908.130 1747.000 908.410 1751.000 ;
    END
  END out_data_flat[233]
  PIN out_data_flat[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 911.350 1747.000 911.630 1751.000 ;
    END
  END out_data_flat[234]
  PIN out_data_flat[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 917.790 1747.000 918.070 1751.000 ;
    END
  END out_data_flat[235]
  PIN out_data_flat[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 901.690 1747.000 901.970 1751.000 ;
    END
  END out_data_flat[236]
  PIN out_data_flat[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 904.910 1747.000 905.190 1751.000 ;
    END
  END out_data_flat[237]
  PIN out_data_flat[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 898.470 1747.000 898.750 1751.000 ;
    END
  END out_data_flat[238]
  PIN out_data_flat[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 895.250 1747.000 895.530 1751.000 ;
    END
  END out_data_flat[239]
  PIN out_data_flat[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 837.290 0.000 837.570 4.000 ;
    END
  END out_data_flat[23]
  PIN out_data_flat[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 836.440 4.000 837.040 ;
    END
  END out_data_flat[240]
  PIN out_data_flat[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 812.640 4.000 813.240 ;
    END
  END out_data_flat[241]
  PIN out_data_flat[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 785.440 4.000 786.040 ;
    END
  END out_data_flat[242]
  PIN out_data_flat[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 751.440 4.000 752.040 ;
    END
  END out_data_flat[243]
  PIN out_data_flat[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 581.440 4.000 582.040 ;
    END
  END out_data_flat[244]
  PIN out_data_flat[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END out_data_flat[245]
  PIN out_data_flat[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 574.640 4.000 575.240 ;
    END
  END out_data_flat[246]
  PIN out_data_flat[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 717.440 4.000 718.040 ;
    END
  END out_data_flat[247]
  PIN out_data_flat[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 921.440 4.000 922.040 ;
    END
  END out_data_flat[248]
  PIN out_data_flat[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 877.240 4.000 877.840 ;
    END
  END out_data_flat[249]
  PIN out_data_flat[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 949.990 1747.000 950.270 1751.000 ;
    END
  END out_data_flat[24]
  PIN out_data_flat[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 938.440 4.000 939.040 ;
    END
  END out_data_flat[250]
  PIN out_data_flat[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 965.640 4.000 966.240 ;
    END
  END out_data_flat[251]
  PIN out_data_flat[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 615.110 1747.000 615.390 1751.000 ;
    END
  END out_data_flat[252]
  PIN out_data_flat[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 624.770 1747.000 625.050 1751.000 ;
    END
  END out_data_flat[253]
  PIN out_data_flat[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 605.450 1747.000 605.730 1751.000 ;
    END
  END out_data_flat[254]
  PIN out_data_flat[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1013.240 4.000 1013.840 ;
    END
  END out_data_flat[255]
  PIN out_data_flat[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 866.270 1747.000 866.550 1751.000 ;
    END
  END out_data_flat[25]
  PIN out_data_flat[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 879.150 1747.000 879.430 1751.000 ;
    END
  END out_data_flat[26]
  PIN out_data_flat[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 869.490 1747.000 869.770 1751.000 ;
    END
  END out_data_flat[27]
  PIN out_data_flat[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 937.110 1747.000 937.390 1751.000 ;
    END
  END out_data_flat[28]
  PIN out_data_flat[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 863.050 1747.000 863.330 1751.000 ;
    END
  END out_data_flat[29]
  PIN out_data_flat[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 816.040 1751.000 816.640 ;
    END
  END out_data_flat[2]
  PIN out_data_flat[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 959.650 1747.000 959.930 1751.000 ;
    END
  END out_data_flat[30]
  PIN out_data_flat[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 814.750 1747.000 815.030 1751.000 ;
    END
  END out_data_flat[31]
  PIN out_data_flat[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 833.040 1751.000 833.640 ;
    END
  END out_data_flat[32]
  PIN out_data_flat[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 829.640 1751.000 830.240 ;
    END
  END out_data_flat[33]
  PIN out_data_flat[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 778.640 1751.000 779.240 ;
    END
  END out_data_flat[34]
  PIN out_data_flat[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 768.440 1751.000 769.040 ;
    END
  END out_data_flat[35]
  PIN out_data_flat[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1136.750 0.000 1137.030 4.000 ;
    END
  END out_data_flat[36]
  PIN out_data_flat[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1123.870 0.000 1124.150 4.000 ;
    END
  END out_data_flat[37]
  PIN out_data_flat[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 717.440 1751.000 718.040 ;
    END
  END out_data_flat[38]
  PIN out_data_flat[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 748.040 1751.000 748.640 ;
    END
  END out_data_flat[39]
  PIN out_data_flat[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 785.440 1751.000 786.040 ;
    END
  END out_data_flat[3]
  PIN out_data_flat[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 822.840 1751.000 823.440 ;
    END
  END out_data_flat[40]
  PIN out_data_flat[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 754.840 1751.000 755.440 ;
    END
  END out_data_flat[41]
  PIN out_data_flat[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 945.240 1751.000 945.840 ;
    END
  END out_data_flat[42]
  PIN out_data_flat[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 996.240 1751.000 996.840 ;
    END
  END out_data_flat[43]
  PIN out_data_flat[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1101.640 1751.000 1102.240 ;
    END
  END out_data_flat[44]
  PIN out_data_flat[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1111.840 1751.000 1112.440 ;
    END
  END out_data_flat[45]
  PIN out_data_flat[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1088.040 1751.000 1088.640 ;
    END
  END out_data_flat[46]
  PIN out_data_flat[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1139.040 1751.000 1139.640 ;
    END
  END out_data_flat[47]
  PIN out_data_flat[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 856.840 4.000 857.440 ;
    END
  END out_data_flat[48]
  PIN out_data_flat[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 826.240 4.000 826.840 ;
    END
  END out_data_flat[49]
  PIN out_data_flat[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1139.970 0.000 1140.250 4.000 ;
    END
  END out_data_flat[4]
  PIN out_data_flat[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 795.640 4.000 796.240 ;
    END
  END out_data_flat[50]
  PIN out_data_flat[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.240 4.000 741.840 ;
    END
  END out_data_flat[51]
  PIN out_data_flat[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 798.650 0.000 798.930 4.000 ;
    END
  END out_data_flat[52]
  PIN out_data_flat[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 801.870 0.000 802.150 4.000 ;
    END
  END out_data_flat[53]
  PIN out_data_flat[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 795.430 0.000 795.710 4.000 ;
    END
  END out_data_flat[54]
  PIN out_data_flat[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 710.640 4.000 711.240 ;
    END
  END out_data_flat[55]
  PIN out_data_flat[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 850.170 1747.000 850.450 1751.000 ;
    END
  END out_data_flat[56]
  PIN out_data_flat[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 801.870 1747.000 802.150 1751.000 ;
    END
  END out_data_flat[57]
  PIN out_data_flat[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 962.870 1747.000 963.150 1751.000 ;
    END
  END out_data_flat[58]
  PIN out_data_flat[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 808.310 1747.000 808.590 1751.000 ;
    END
  END out_data_flat[59]
  PIN out_data_flat[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 724.240 1751.000 724.840 ;
    END
  END out_data_flat[5]
  PIN out_data_flat[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 846.950 1747.000 847.230 1751.000 ;
    END
  END out_data_flat[60]
  PIN out_data_flat[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 805.090 1747.000 805.370 1751.000 ;
    END
  END out_data_flat[61]
  PIN out_data_flat[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 811.530 1747.000 811.810 1751.000 ;
    END
  END out_data_flat[62]
  PIN out_data_flat[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 792.210 1747.000 792.490 1751.000 ;
    END
  END out_data_flat[63]
  PIN out_data_flat[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 863.640 1751.000 864.240 ;
    END
  END out_data_flat[64]
  PIN out_data_flat[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 836.440 1751.000 837.040 ;
    END
  END out_data_flat[65]
  PIN out_data_flat[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 788.840 1751.000 789.440 ;
    END
  END out_data_flat[66]
  PIN out_data_flat[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 775.240 1751.000 775.840 ;
    END
  END out_data_flat[67]
  PIN out_data_flat[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1110.990 0.000 1111.270 4.000 ;
    END
  END out_data_flat[68]
  PIN out_data_flat[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1107.770 0.000 1108.050 4.000 ;
    END
  END out_data_flat[69]
  PIN out_data_flat[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 731.040 1751.000 731.640 ;
    END
  END out_data_flat[6]
  PIN out_data_flat[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1117.430 0.000 1117.710 4.000 ;
    END
  END out_data_flat[70]
  PIN out_data_flat[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1114.210 0.000 1114.490 4.000 ;
    END
  END out_data_flat[71]
  PIN out_data_flat[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 873.840 1751.000 874.440 ;
    END
  END out_data_flat[72]
  PIN out_data_flat[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 734.440 1751.000 735.040 ;
    END
  END out_data_flat[73]
  PIN out_data_flat[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 982.640 1751.000 983.240 ;
    END
  END out_data_flat[74]
  PIN out_data_flat[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1071.040 1751.000 1071.640 ;
    END
  END out_data_flat[75]
  PIN out_data_flat[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1162.840 1751.000 1163.440 ;
    END
  END out_data_flat[76]
  PIN out_data_flat[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1108.440 1751.000 1109.040 ;
    END
  END out_data_flat[77]
  PIN out_data_flat[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1098.240 1751.000 1098.840 ;
    END
  END out_data_flat[78]
  PIN out_data_flat[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 1050.640 1751.000 1051.240 ;
    END
  END out_data_flat[79]
  PIN out_data_flat[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 758.240 1751.000 758.840 ;
    END
  END out_data_flat[7]
  PIN out_data_flat[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 867.040 4.000 867.640 ;
    END
  END out_data_flat[80]
  PIN out_data_flat[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 822.840 4.000 823.440 ;
    END
  END out_data_flat[81]
  PIN out_data_flat[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.240 4.000 792.840 ;
    END
  END out_data_flat[82]
  PIN out_data_flat[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.840 4.000 704.440 ;
    END
  END out_data_flat[83]
  PIN out_data_flat[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END out_data_flat[84]
  PIN out_data_flat[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END out_data_flat[85]
  PIN out_data_flat[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 642.640 4.000 643.240 ;
    END
  END out_data_flat[86]
  PIN out_data_flat[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 700.440 4.000 701.040 ;
    END
  END out_data_flat[87]
  PIN out_data_flat[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 766.450 1747.000 766.730 1751.000 ;
    END
  END out_data_flat[88]
  PIN out_data_flat[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 795.430 1747.000 795.710 1751.000 ;
    END
  END out_data_flat[89]
  PIN out_data_flat[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 799.040 1751.000 799.640 ;
    END
  END out_data_flat[8]
  PIN out_data_flat[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 731.030 1747.000 731.310 1751.000 ;
    END
  END out_data_flat[90]
  PIN out_data_flat[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 740.690 1747.000 740.970 1751.000 ;
    END
  END out_data_flat[91]
  PIN out_data_flat[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 760.010 1747.000 760.290 1751.000 ;
    END
  END out_data_flat[92]
  PIN out_data_flat[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 756.790 1747.000 757.070 1751.000 ;
    END
  END out_data_flat[93]
  PIN out_data_flat[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 763.230 1747.000 763.510 1751.000 ;
    END
  END out_data_flat[94]
  PIN out_data_flat[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 750.350 1747.000 750.630 1751.000 ;
    END
  END out_data_flat[95]
  PIN out_data_flat[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 802.440 1751.000 803.040 ;
    END
  END out_data_flat[96]
  PIN out_data_flat[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 812.640 1751.000 813.240 ;
    END
  END out_data_flat[97]
  PIN out_data_flat[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1069.130 0.000 1069.410 4.000 ;
    END
  END out_data_flat[98]
  PIN out_data_flat[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1065.910 0.000 1066.190 4.000 ;
    END
  END out_data_flat[99]
  PIN out_data_flat[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1747.000 907.840 1751.000 908.440 ;
    END
  END out_data_flat[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1060.840 4.000 1061.440 ;
    END
  END rst
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 1745.430 1738.270 ;
      LAYER li1 ;
        RECT 5.520 10.795 1745.240 1738.165 ;
      LAYER met1 ;
        RECT 4.210 9.220 1745.240 1738.320 ;
      LAYER met2 ;
        RECT 4.230 1746.720 595.510 1747.330 ;
        RECT 596.350 1746.720 605.170 1747.330 ;
        RECT 606.010 1746.720 608.390 1747.330 ;
        RECT 609.230 1746.720 611.610 1747.330 ;
        RECT 612.450 1746.720 614.830 1747.330 ;
        RECT 615.670 1746.720 618.050 1747.330 ;
        RECT 618.890 1746.720 621.270 1747.330 ;
        RECT 622.110 1746.720 624.490 1747.330 ;
        RECT 625.330 1746.720 627.710 1747.330 ;
        RECT 628.550 1746.720 630.930 1747.330 ;
        RECT 631.770 1746.720 634.150 1747.330 ;
        RECT 634.990 1746.720 637.370 1747.330 ;
        RECT 638.210 1746.720 640.590 1747.330 ;
        RECT 641.430 1746.720 643.810 1747.330 ;
        RECT 644.650 1746.720 647.030 1747.330 ;
        RECT 647.870 1746.720 650.250 1747.330 ;
        RECT 651.090 1746.720 653.470 1747.330 ;
        RECT 654.310 1746.720 656.690 1747.330 ;
        RECT 657.530 1746.720 659.910 1747.330 ;
        RECT 660.750 1746.720 663.130 1747.330 ;
        RECT 663.970 1746.720 666.350 1747.330 ;
        RECT 667.190 1746.720 669.570 1747.330 ;
        RECT 670.410 1746.720 672.790 1747.330 ;
        RECT 673.630 1746.720 676.010 1747.330 ;
        RECT 676.850 1746.720 679.230 1747.330 ;
        RECT 680.070 1746.720 682.450 1747.330 ;
        RECT 683.290 1746.720 685.670 1747.330 ;
        RECT 686.510 1746.720 688.890 1747.330 ;
        RECT 689.730 1746.720 692.110 1747.330 ;
        RECT 692.950 1746.720 695.330 1747.330 ;
        RECT 696.170 1746.720 698.550 1747.330 ;
        RECT 699.390 1746.720 701.770 1747.330 ;
        RECT 702.610 1746.720 704.990 1747.330 ;
        RECT 705.830 1746.720 708.210 1747.330 ;
        RECT 709.050 1746.720 711.430 1747.330 ;
        RECT 712.270 1746.720 714.650 1747.330 ;
        RECT 715.490 1746.720 717.870 1747.330 ;
        RECT 718.710 1746.720 721.090 1747.330 ;
        RECT 721.930 1746.720 724.310 1747.330 ;
        RECT 725.150 1746.720 727.530 1747.330 ;
        RECT 728.370 1746.720 730.750 1747.330 ;
        RECT 731.590 1746.720 733.970 1747.330 ;
        RECT 734.810 1746.720 737.190 1747.330 ;
        RECT 738.030 1746.720 740.410 1747.330 ;
        RECT 741.250 1746.720 743.630 1747.330 ;
        RECT 744.470 1746.720 746.850 1747.330 ;
        RECT 747.690 1746.720 750.070 1747.330 ;
        RECT 750.910 1746.720 753.290 1747.330 ;
        RECT 754.130 1746.720 756.510 1747.330 ;
        RECT 757.350 1746.720 759.730 1747.330 ;
        RECT 760.570 1746.720 762.950 1747.330 ;
        RECT 763.790 1746.720 766.170 1747.330 ;
        RECT 767.010 1746.720 769.390 1747.330 ;
        RECT 770.230 1746.720 772.610 1747.330 ;
        RECT 773.450 1746.720 775.830 1747.330 ;
        RECT 776.670 1746.720 779.050 1747.330 ;
        RECT 779.890 1746.720 782.270 1747.330 ;
        RECT 783.110 1746.720 785.490 1747.330 ;
        RECT 786.330 1746.720 788.710 1747.330 ;
        RECT 789.550 1746.720 791.930 1747.330 ;
        RECT 792.770 1746.720 795.150 1747.330 ;
        RECT 795.990 1746.720 798.370 1747.330 ;
        RECT 799.210 1746.720 801.590 1747.330 ;
        RECT 802.430 1746.720 804.810 1747.330 ;
        RECT 805.650 1746.720 808.030 1747.330 ;
        RECT 808.870 1746.720 811.250 1747.330 ;
        RECT 812.090 1746.720 814.470 1747.330 ;
        RECT 815.310 1746.720 817.690 1747.330 ;
        RECT 818.530 1746.720 820.910 1747.330 ;
        RECT 821.750 1746.720 824.130 1747.330 ;
        RECT 824.970 1746.720 827.350 1747.330 ;
        RECT 828.190 1746.720 830.570 1747.330 ;
        RECT 831.410 1746.720 833.790 1747.330 ;
        RECT 834.630 1746.720 837.010 1747.330 ;
        RECT 837.850 1746.720 840.230 1747.330 ;
        RECT 841.070 1746.720 843.450 1747.330 ;
        RECT 844.290 1746.720 846.670 1747.330 ;
        RECT 847.510 1746.720 849.890 1747.330 ;
        RECT 850.730 1746.720 853.110 1747.330 ;
        RECT 853.950 1746.720 856.330 1747.330 ;
        RECT 857.170 1746.720 859.550 1747.330 ;
        RECT 860.390 1746.720 862.770 1747.330 ;
        RECT 863.610 1746.720 865.990 1747.330 ;
        RECT 866.830 1746.720 869.210 1747.330 ;
        RECT 870.050 1746.720 872.430 1747.330 ;
        RECT 873.270 1746.720 875.650 1747.330 ;
        RECT 876.490 1746.720 878.870 1747.330 ;
        RECT 879.710 1746.720 882.090 1747.330 ;
        RECT 882.930 1746.720 885.310 1747.330 ;
        RECT 886.150 1746.720 888.530 1747.330 ;
        RECT 889.370 1746.720 891.750 1747.330 ;
        RECT 892.590 1746.720 894.970 1747.330 ;
        RECT 895.810 1746.720 898.190 1747.330 ;
        RECT 899.030 1746.720 901.410 1747.330 ;
        RECT 902.250 1746.720 904.630 1747.330 ;
        RECT 905.470 1746.720 907.850 1747.330 ;
        RECT 908.690 1746.720 911.070 1747.330 ;
        RECT 911.910 1746.720 914.290 1747.330 ;
        RECT 915.130 1746.720 917.510 1747.330 ;
        RECT 918.350 1746.720 920.730 1747.330 ;
        RECT 921.570 1746.720 923.950 1747.330 ;
        RECT 924.790 1746.720 927.170 1747.330 ;
        RECT 928.010 1746.720 930.390 1747.330 ;
        RECT 931.230 1746.720 933.610 1747.330 ;
        RECT 934.450 1746.720 936.830 1747.330 ;
        RECT 937.670 1746.720 940.050 1747.330 ;
        RECT 940.890 1746.720 943.270 1747.330 ;
        RECT 944.110 1746.720 946.490 1747.330 ;
        RECT 947.330 1746.720 949.710 1747.330 ;
        RECT 950.550 1746.720 952.930 1747.330 ;
        RECT 953.770 1746.720 956.150 1747.330 ;
        RECT 956.990 1746.720 959.370 1747.330 ;
        RECT 960.210 1746.720 962.590 1747.330 ;
        RECT 963.430 1746.720 965.810 1747.330 ;
        RECT 966.650 1746.720 969.030 1747.330 ;
        RECT 969.870 1746.720 994.790 1747.330 ;
        RECT 995.630 1746.720 1743.770 1747.330 ;
        RECT 4.230 4.280 1743.770 1746.720 ;
        RECT 4.230 4.000 759.730 4.280 ;
        RECT 760.570 4.000 762.950 4.280 ;
        RECT 763.790 4.000 766.170 4.280 ;
        RECT 767.010 4.000 769.390 4.280 ;
        RECT 770.230 4.000 772.610 4.280 ;
        RECT 773.450 4.000 775.830 4.280 ;
        RECT 776.670 4.000 779.050 4.280 ;
        RECT 779.890 4.000 782.270 4.280 ;
        RECT 783.110 4.000 785.490 4.280 ;
        RECT 786.330 4.000 788.710 4.280 ;
        RECT 789.550 4.000 791.930 4.280 ;
        RECT 792.770 4.000 795.150 4.280 ;
        RECT 795.990 4.000 798.370 4.280 ;
        RECT 799.210 4.000 801.590 4.280 ;
        RECT 802.430 4.000 804.810 4.280 ;
        RECT 805.650 4.000 808.030 4.280 ;
        RECT 808.870 4.000 811.250 4.280 ;
        RECT 812.090 4.000 814.470 4.280 ;
        RECT 815.310 4.000 817.690 4.280 ;
        RECT 818.530 4.000 820.910 4.280 ;
        RECT 821.750 4.000 824.130 4.280 ;
        RECT 824.970 4.000 827.350 4.280 ;
        RECT 828.190 4.000 830.570 4.280 ;
        RECT 831.410 4.000 833.790 4.280 ;
        RECT 834.630 4.000 837.010 4.280 ;
        RECT 837.850 4.000 840.230 4.280 ;
        RECT 841.070 4.000 843.450 4.280 ;
        RECT 844.290 4.000 846.670 4.280 ;
        RECT 847.510 4.000 849.890 4.280 ;
        RECT 850.730 4.000 853.110 4.280 ;
        RECT 853.950 4.000 856.330 4.280 ;
        RECT 857.170 4.000 859.550 4.280 ;
        RECT 860.390 4.000 862.770 4.280 ;
        RECT 863.610 4.000 865.990 4.280 ;
        RECT 866.830 4.000 869.210 4.280 ;
        RECT 870.050 4.000 872.430 4.280 ;
        RECT 873.270 4.000 875.650 4.280 ;
        RECT 876.490 4.000 878.870 4.280 ;
        RECT 879.710 4.000 882.090 4.280 ;
        RECT 882.930 4.000 885.310 4.280 ;
        RECT 886.150 4.000 888.530 4.280 ;
        RECT 889.370 4.000 891.750 4.280 ;
        RECT 892.590 4.000 894.970 4.280 ;
        RECT 895.810 4.000 898.190 4.280 ;
        RECT 899.030 4.000 901.410 4.280 ;
        RECT 902.250 4.000 904.630 4.280 ;
        RECT 905.470 4.000 907.850 4.280 ;
        RECT 908.690 4.000 911.070 4.280 ;
        RECT 911.910 4.000 914.290 4.280 ;
        RECT 915.130 4.000 917.510 4.280 ;
        RECT 918.350 4.000 920.730 4.280 ;
        RECT 921.570 4.000 923.950 4.280 ;
        RECT 924.790 4.000 927.170 4.280 ;
        RECT 928.010 4.000 930.390 4.280 ;
        RECT 931.230 4.000 933.610 4.280 ;
        RECT 934.450 4.000 936.830 4.280 ;
        RECT 937.670 4.000 940.050 4.280 ;
        RECT 940.890 4.000 943.270 4.280 ;
        RECT 944.110 4.000 946.490 4.280 ;
        RECT 947.330 4.000 949.710 4.280 ;
        RECT 950.550 4.000 952.930 4.280 ;
        RECT 953.770 4.000 956.150 4.280 ;
        RECT 956.990 4.000 959.370 4.280 ;
        RECT 960.210 4.000 962.590 4.280 ;
        RECT 963.430 4.000 965.810 4.280 ;
        RECT 966.650 4.000 969.030 4.280 ;
        RECT 969.870 4.000 972.250 4.280 ;
        RECT 973.090 4.000 975.470 4.280 ;
        RECT 976.310 4.000 978.690 4.280 ;
        RECT 979.530 4.000 981.910 4.280 ;
        RECT 982.750 4.000 985.130 4.280 ;
        RECT 985.970 4.000 988.350 4.280 ;
        RECT 989.190 4.000 991.570 4.280 ;
        RECT 992.410 4.000 994.790 4.280 ;
        RECT 995.630 4.000 998.010 4.280 ;
        RECT 998.850 4.000 1001.230 4.280 ;
        RECT 1002.070 4.000 1004.450 4.280 ;
        RECT 1005.290 4.000 1007.670 4.280 ;
        RECT 1008.510 4.000 1010.890 4.280 ;
        RECT 1011.730 4.000 1014.110 4.280 ;
        RECT 1014.950 4.000 1017.330 4.280 ;
        RECT 1018.170 4.000 1020.550 4.280 ;
        RECT 1021.390 4.000 1023.770 4.280 ;
        RECT 1024.610 4.000 1026.990 4.280 ;
        RECT 1027.830 4.000 1030.210 4.280 ;
        RECT 1031.050 4.000 1033.430 4.280 ;
        RECT 1034.270 4.000 1036.650 4.280 ;
        RECT 1037.490 4.000 1039.870 4.280 ;
        RECT 1040.710 4.000 1043.090 4.280 ;
        RECT 1043.930 4.000 1046.310 4.280 ;
        RECT 1047.150 4.000 1049.530 4.280 ;
        RECT 1050.370 4.000 1052.750 4.280 ;
        RECT 1053.590 4.000 1055.970 4.280 ;
        RECT 1056.810 4.000 1059.190 4.280 ;
        RECT 1060.030 4.000 1062.410 4.280 ;
        RECT 1063.250 4.000 1065.630 4.280 ;
        RECT 1066.470 4.000 1068.850 4.280 ;
        RECT 1069.690 4.000 1072.070 4.280 ;
        RECT 1072.910 4.000 1075.290 4.280 ;
        RECT 1076.130 4.000 1078.510 4.280 ;
        RECT 1079.350 4.000 1081.730 4.280 ;
        RECT 1082.570 4.000 1084.950 4.280 ;
        RECT 1085.790 4.000 1088.170 4.280 ;
        RECT 1089.010 4.000 1091.390 4.280 ;
        RECT 1092.230 4.000 1094.610 4.280 ;
        RECT 1095.450 4.000 1097.830 4.280 ;
        RECT 1098.670 4.000 1101.050 4.280 ;
        RECT 1101.890 4.000 1104.270 4.280 ;
        RECT 1105.110 4.000 1107.490 4.280 ;
        RECT 1108.330 4.000 1110.710 4.280 ;
        RECT 1111.550 4.000 1113.930 4.280 ;
        RECT 1114.770 4.000 1117.150 4.280 ;
        RECT 1117.990 4.000 1120.370 4.280 ;
        RECT 1121.210 4.000 1123.590 4.280 ;
        RECT 1124.430 4.000 1126.810 4.280 ;
        RECT 1127.650 4.000 1130.030 4.280 ;
        RECT 1130.870 4.000 1133.250 4.280 ;
        RECT 1134.090 4.000 1136.470 4.280 ;
        RECT 1137.310 4.000 1139.690 4.280 ;
        RECT 1140.530 4.000 1152.570 4.280 ;
        RECT 1153.410 4.000 1743.770 4.280 ;
      LAYER met3 ;
        RECT 3.750 1184.240 1747.000 1738.245 ;
        RECT 3.750 1182.840 1746.600 1184.240 ;
        RECT 3.750 1180.840 1747.000 1182.840 ;
        RECT 3.750 1179.440 1746.600 1180.840 ;
        RECT 3.750 1177.440 1747.000 1179.440 ;
        RECT 3.750 1176.040 1746.600 1177.440 ;
        RECT 3.750 1174.040 1747.000 1176.040 ;
        RECT 3.750 1172.640 1746.600 1174.040 ;
        RECT 3.750 1170.640 1747.000 1172.640 ;
        RECT 3.750 1169.240 1746.600 1170.640 ;
        RECT 3.750 1167.240 1747.000 1169.240 ;
        RECT 3.750 1165.840 1746.600 1167.240 ;
        RECT 3.750 1163.840 1747.000 1165.840 ;
        RECT 3.750 1162.440 1746.600 1163.840 ;
        RECT 3.750 1160.440 1747.000 1162.440 ;
        RECT 3.750 1159.040 1746.600 1160.440 ;
        RECT 3.750 1157.040 1747.000 1159.040 ;
        RECT 3.750 1155.640 1746.600 1157.040 ;
        RECT 3.750 1153.640 1747.000 1155.640 ;
        RECT 3.750 1152.240 1746.600 1153.640 ;
        RECT 3.750 1150.240 1747.000 1152.240 ;
        RECT 3.750 1148.840 1746.600 1150.240 ;
        RECT 3.750 1146.840 1747.000 1148.840 ;
        RECT 3.750 1145.440 1746.600 1146.840 ;
        RECT 3.750 1143.440 1747.000 1145.440 ;
        RECT 3.750 1142.040 1746.600 1143.440 ;
        RECT 3.750 1140.040 1747.000 1142.040 ;
        RECT 3.750 1138.640 1746.600 1140.040 ;
        RECT 3.750 1136.640 1747.000 1138.640 ;
        RECT 3.750 1135.240 1746.600 1136.640 ;
        RECT 3.750 1133.240 1747.000 1135.240 ;
        RECT 3.750 1131.840 1746.600 1133.240 ;
        RECT 3.750 1129.840 1747.000 1131.840 ;
        RECT 3.750 1128.440 1746.600 1129.840 ;
        RECT 3.750 1126.440 1747.000 1128.440 ;
        RECT 3.750 1125.040 1746.600 1126.440 ;
        RECT 3.750 1123.040 1747.000 1125.040 ;
        RECT 3.750 1121.640 1746.600 1123.040 ;
        RECT 3.750 1119.640 1747.000 1121.640 ;
        RECT 3.750 1118.240 1746.600 1119.640 ;
        RECT 3.750 1116.240 1747.000 1118.240 ;
        RECT 3.750 1114.840 1746.600 1116.240 ;
        RECT 3.750 1112.840 1747.000 1114.840 ;
        RECT 3.750 1111.440 1746.600 1112.840 ;
        RECT 3.750 1109.440 1747.000 1111.440 ;
        RECT 3.750 1108.040 1746.600 1109.440 ;
        RECT 3.750 1106.040 1747.000 1108.040 ;
        RECT 3.750 1104.640 1746.600 1106.040 ;
        RECT 3.750 1102.640 1747.000 1104.640 ;
        RECT 3.750 1101.240 1746.600 1102.640 ;
        RECT 3.750 1099.240 1747.000 1101.240 ;
        RECT 3.750 1097.840 1746.600 1099.240 ;
        RECT 3.750 1095.840 1747.000 1097.840 ;
        RECT 3.750 1094.440 1746.600 1095.840 ;
        RECT 3.750 1092.440 1747.000 1094.440 ;
        RECT 3.750 1091.040 1746.600 1092.440 ;
        RECT 3.750 1089.040 1747.000 1091.040 ;
        RECT 3.750 1087.640 1746.600 1089.040 ;
        RECT 3.750 1085.640 1747.000 1087.640 ;
        RECT 3.750 1084.240 1746.600 1085.640 ;
        RECT 3.750 1082.240 1747.000 1084.240 ;
        RECT 3.750 1080.840 1746.600 1082.240 ;
        RECT 3.750 1078.840 1747.000 1080.840 ;
        RECT 3.750 1077.440 1746.600 1078.840 ;
        RECT 3.750 1075.440 1747.000 1077.440 ;
        RECT 3.750 1074.040 1746.600 1075.440 ;
        RECT 3.750 1072.040 1747.000 1074.040 ;
        RECT 3.750 1070.640 1746.600 1072.040 ;
        RECT 3.750 1068.640 1747.000 1070.640 ;
        RECT 4.400 1067.240 1746.600 1068.640 ;
        RECT 3.750 1065.240 1747.000 1067.240 ;
        RECT 4.400 1063.840 1746.600 1065.240 ;
        RECT 3.750 1061.840 1747.000 1063.840 ;
        RECT 4.400 1060.440 1746.600 1061.840 ;
        RECT 3.750 1058.440 1747.000 1060.440 ;
        RECT 3.750 1057.040 1746.600 1058.440 ;
        RECT 3.750 1055.040 1747.000 1057.040 ;
        RECT 3.750 1053.640 1746.600 1055.040 ;
        RECT 3.750 1051.640 1747.000 1053.640 ;
        RECT 3.750 1050.240 1746.600 1051.640 ;
        RECT 3.750 1048.240 1747.000 1050.240 ;
        RECT 3.750 1046.840 1746.600 1048.240 ;
        RECT 3.750 1044.840 1747.000 1046.840 ;
        RECT 3.750 1043.440 1746.600 1044.840 ;
        RECT 3.750 1041.440 1747.000 1043.440 ;
        RECT 3.750 1040.040 1746.600 1041.440 ;
        RECT 3.750 1038.040 1747.000 1040.040 ;
        RECT 3.750 1036.640 1746.600 1038.040 ;
        RECT 3.750 1034.640 1747.000 1036.640 ;
        RECT 3.750 1033.240 1746.600 1034.640 ;
        RECT 3.750 1031.240 1747.000 1033.240 ;
        RECT 3.750 1029.840 1746.600 1031.240 ;
        RECT 3.750 1027.840 1747.000 1029.840 ;
        RECT 3.750 1026.440 1746.600 1027.840 ;
        RECT 3.750 1024.440 1747.000 1026.440 ;
        RECT 3.750 1023.040 1746.600 1024.440 ;
        RECT 3.750 1021.040 1747.000 1023.040 ;
        RECT 4.400 1019.640 1746.600 1021.040 ;
        RECT 3.750 1017.640 1747.000 1019.640 ;
        RECT 3.750 1016.240 1746.600 1017.640 ;
        RECT 3.750 1014.240 1747.000 1016.240 ;
        RECT 4.400 1012.840 1746.600 1014.240 ;
        RECT 3.750 1010.840 1747.000 1012.840 ;
        RECT 4.400 1009.440 1746.600 1010.840 ;
        RECT 3.750 1007.440 1747.000 1009.440 ;
        RECT 4.400 1006.040 1746.600 1007.440 ;
        RECT 3.750 1004.040 1747.000 1006.040 ;
        RECT 4.400 1002.640 1746.600 1004.040 ;
        RECT 3.750 1000.640 1747.000 1002.640 ;
        RECT 4.400 999.240 1746.600 1000.640 ;
        RECT 3.750 997.240 1747.000 999.240 ;
        RECT 4.400 995.840 1746.600 997.240 ;
        RECT 3.750 993.840 1747.000 995.840 ;
        RECT 4.400 992.440 1746.600 993.840 ;
        RECT 3.750 990.440 1747.000 992.440 ;
        RECT 4.400 989.040 1746.600 990.440 ;
        RECT 3.750 987.040 1747.000 989.040 ;
        RECT 4.400 985.640 1746.600 987.040 ;
        RECT 3.750 983.640 1747.000 985.640 ;
        RECT 4.400 982.240 1746.600 983.640 ;
        RECT 3.750 980.240 1747.000 982.240 ;
        RECT 4.400 978.840 1746.600 980.240 ;
        RECT 3.750 976.840 1747.000 978.840 ;
        RECT 4.400 975.440 1746.600 976.840 ;
        RECT 3.750 973.440 1747.000 975.440 ;
        RECT 4.400 972.040 1746.600 973.440 ;
        RECT 3.750 970.040 1747.000 972.040 ;
        RECT 4.400 968.640 1746.600 970.040 ;
        RECT 3.750 966.640 1747.000 968.640 ;
        RECT 4.400 965.240 1746.600 966.640 ;
        RECT 3.750 963.240 1747.000 965.240 ;
        RECT 4.400 961.840 1746.600 963.240 ;
        RECT 3.750 959.840 1747.000 961.840 ;
        RECT 4.400 958.440 1746.600 959.840 ;
        RECT 3.750 956.440 1747.000 958.440 ;
        RECT 4.400 955.040 1746.600 956.440 ;
        RECT 3.750 953.040 1747.000 955.040 ;
        RECT 4.400 951.640 1746.600 953.040 ;
        RECT 3.750 949.640 1747.000 951.640 ;
        RECT 4.400 948.240 1746.600 949.640 ;
        RECT 3.750 946.240 1747.000 948.240 ;
        RECT 4.400 944.840 1746.600 946.240 ;
        RECT 3.750 942.840 1747.000 944.840 ;
        RECT 4.400 941.440 1746.600 942.840 ;
        RECT 3.750 939.440 1747.000 941.440 ;
        RECT 4.400 938.040 1746.600 939.440 ;
        RECT 3.750 936.040 1747.000 938.040 ;
        RECT 4.400 934.640 1746.600 936.040 ;
        RECT 3.750 932.640 1747.000 934.640 ;
        RECT 4.400 931.240 1746.600 932.640 ;
        RECT 3.750 929.240 1747.000 931.240 ;
        RECT 4.400 927.840 1746.600 929.240 ;
        RECT 3.750 925.840 1747.000 927.840 ;
        RECT 4.400 924.440 1746.600 925.840 ;
        RECT 3.750 922.440 1747.000 924.440 ;
        RECT 4.400 921.040 1746.600 922.440 ;
        RECT 3.750 919.040 1747.000 921.040 ;
        RECT 4.400 917.640 1746.600 919.040 ;
        RECT 3.750 915.640 1747.000 917.640 ;
        RECT 4.400 914.240 1746.600 915.640 ;
        RECT 3.750 912.240 1747.000 914.240 ;
        RECT 4.400 910.840 1746.600 912.240 ;
        RECT 3.750 908.840 1747.000 910.840 ;
        RECT 4.400 907.440 1746.600 908.840 ;
        RECT 3.750 905.440 1747.000 907.440 ;
        RECT 4.400 904.040 1746.600 905.440 ;
        RECT 3.750 902.040 1747.000 904.040 ;
        RECT 4.400 900.640 1746.600 902.040 ;
        RECT 3.750 898.640 1747.000 900.640 ;
        RECT 4.400 897.240 1746.600 898.640 ;
        RECT 3.750 895.240 1747.000 897.240 ;
        RECT 4.400 893.840 1746.600 895.240 ;
        RECT 3.750 891.840 1747.000 893.840 ;
        RECT 4.400 890.440 1746.600 891.840 ;
        RECT 3.750 888.440 1747.000 890.440 ;
        RECT 4.400 887.040 1746.600 888.440 ;
        RECT 3.750 885.040 1747.000 887.040 ;
        RECT 4.400 883.640 1746.600 885.040 ;
        RECT 3.750 881.640 1747.000 883.640 ;
        RECT 4.400 880.240 1746.600 881.640 ;
        RECT 3.750 878.240 1747.000 880.240 ;
        RECT 4.400 876.840 1746.600 878.240 ;
        RECT 3.750 874.840 1747.000 876.840 ;
        RECT 4.400 873.440 1746.600 874.840 ;
        RECT 3.750 871.440 1747.000 873.440 ;
        RECT 4.400 870.040 1746.600 871.440 ;
        RECT 3.750 868.040 1747.000 870.040 ;
        RECT 4.400 866.640 1746.600 868.040 ;
        RECT 3.750 864.640 1747.000 866.640 ;
        RECT 4.400 863.240 1746.600 864.640 ;
        RECT 3.750 861.240 1747.000 863.240 ;
        RECT 4.400 859.840 1746.600 861.240 ;
        RECT 3.750 857.840 1747.000 859.840 ;
        RECT 4.400 856.440 1746.600 857.840 ;
        RECT 3.750 854.440 1747.000 856.440 ;
        RECT 4.400 853.040 1746.600 854.440 ;
        RECT 3.750 851.040 1747.000 853.040 ;
        RECT 4.400 849.640 1746.600 851.040 ;
        RECT 3.750 847.640 1747.000 849.640 ;
        RECT 4.400 846.240 1746.600 847.640 ;
        RECT 3.750 844.240 1747.000 846.240 ;
        RECT 4.400 842.840 1746.600 844.240 ;
        RECT 3.750 840.840 1747.000 842.840 ;
        RECT 4.400 839.440 1746.600 840.840 ;
        RECT 3.750 837.440 1747.000 839.440 ;
        RECT 4.400 836.040 1746.600 837.440 ;
        RECT 3.750 834.040 1747.000 836.040 ;
        RECT 4.400 832.640 1746.600 834.040 ;
        RECT 3.750 830.640 1747.000 832.640 ;
        RECT 4.400 829.240 1746.600 830.640 ;
        RECT 3.750 827.240 1747.000 829.240 ;
        RECT 4.400 825.840 1746.600 827.240 ;
        RECT 3.750 823.840 1747.000 825.840 ;
        RECT 4.400 822.440 1746.600 823.840 ;
        RECT 3.750 820.440 1747.000 822.440 ;
        RECT 4.400 819.040 1746.600 820.440 ;
        RECT 3.750 817.040 1747.000 819.040 ;
        RECT 4.400 815.640 1746.600 817.040 ;
        RECT 3.750 813.640 1747.000 815.640 ;
        RECT 4.400 812.240 1746.600 813.640 ;
        RECT 3.750 810.240 1747.000 812.240 ;
        RECT 4.400 808.840 1746.600 810.240 ;
        RECT 3.750 806.840 1747.000 808.840 ;
        RECT 4.400 805.440 1746.600 806.840 ;
        RECT 3.750 803.440 1747.000 805.440 ;
        RECT 4.400 802.040 1746.600 803.440 ;
        RECT 3.750 800.040 1747.000 802.040 ;
        RECT 4.400 798.640 1746.600 800.040 ;
        RECT 3.750 796.640 1747.000 798.640 ;
        RECT 4.400 795.240 1746.600 796.640 ;
        RECT 3.750 793.240 1747.000 795.240 ;
        RECT 4.400 791.840 1746.600 793.240 ;
        RECT 3.750 789.840 1747.000 791.840 ;
        RECT 4.400 788.440 1746.600 789.840 ;
        RECT 3.750 786.440 1747.000 788.440 ;
        RECT 4.400 785.040 1746.600 786.440 ;
        RECT 3.750 783.040 1747.000 785.040 ;
        RECT 4.400 781.640 1746.600 783.040 ;
        RECT 3.750 779.640 1747.000 781.640 ;
        RECT 4.400 778.240 1746.600 779.640 ;
        RECT 3.750 776.240 1747.000 778.240 ;
        RECT 4.400 774.840 1746.600 776.240 ;
        RECT 3.750 772.840 1747.000 774.840 ;
        RECT 4.400 771.440 1746.600 772.840 ;
        RECT 3.750 769.440 1747.000 771.440 ;
        RECT 4.400 768.040 1746.600 769.440 ;
        RECT 3.750 766.040 1747.000 768.040 ;
        RECT 4.400 764.640 1746.600 766.040 ;
        RECT 3.750 762.640 1747.000 764.640 ;
        RECT 4.400 761.240 1746.600 762.640 ;
        RECT 3.750 759.240 1747.000 761.240 ;
        RECT 4.400 757.840 1746.600 759.240 ;
        RECT 3.750 755.840 1747.000 757.840 ;
        RECT 4.400 754.440 1746.600 755.840 ;
        RECT 3.750 752.440 1747.000 754.440 ;
        RECT 4.400 751.040 1746.600 752.440 ;
        RECT 3.750 749.040 1747.000 751.040 ;
        RECT 4.400 747.640 1746.600 749.040 ;
        RECT 3.750 745.640 1747.000 747.640 ;
        RECT 4.400 744.240 1746.600 745.640 ;
        RECT 3.750 742.240 1747.000 744.240 ;
        RECT 4.400 740.840 1746.600 742.240 ;
        RECT 3.750 738.840 1747.000 740.840 ;
        RECT 4.400 737.440 1746.600 738.840 ;
        RECT 3.750 735.440 1747.000 737.440 ;
        RECT 4.400 734.040 1746.600 735.440 ;
        RECT 3.750 732.040 1747.000 734.040 ;
        RECT 4.400 730.640 1746.600 732.040 ;
        RECT 3.750 728.640 1747.000 730.640 ;
        RECT 4.400 727.240 1747.000 728.640 ;
        RECT 3.750 725.240 1747.000 727.240 ;
        RECT 4.400 723.840 1746.600 725.240 ;
        RECT 3.750 721.840 1747.000 723.840 ;
        RECT 4.400 720.440 1746.600 721.840 ;
        RECT 3.750 718.440 1747.000 720.440 ;
        RECT 4.400 717.040 1746.600 718.440 ;
        RECT 3.750 715.040 1747.000 717.040 ;
        RECT 4.400 713.640 1747.000 715.040 ;
        RECT 3.750 711.640 1747.000 713.640 ;
        RECT 4.400 710.240 1747.000 711.640 ;
        RECT 3.750 708.240 1747.000 710.240 ;
        RECT 4.400 706.840 1747.000 708.240 ;
        RECT 3.750 704.840 1747.000 706.840 ;
        RECT 4.400 703.440 1747.000 704.840 ;
        RECT 3.750 701.440 1747.000 703.440 ;
        RECT 4.400 700.040 1747.000 701.440 ;
        RECT 3.750 698.040 1747.000 700.040 ;
        RECT 4.400 696.640 1747.000 698.040 ;
        RECT 3.750 694.640 1747.000 696.640 ;
        RECT 4.400 693.240 1747.000 694.640 ;
        RECT 3.750 691.240 1747.000 693.240 ;
        RECT 4.400 689.840 1747.000 691.240 ;
        RECT 3.750 687.840 1747.000 689.840 ;
        RECT 4.400 686.440 1747.000 687.840 ;
        RECT 3.750 684.440 1747.000 686.440 ;
        RECT 4.400 683.040 1747.000 684.440 ;
        RECT 3.750 681.040 1747.000 683.040 ;
        RECT 4.400 679.640 1747.000 681.040 ;
        RECT 3.750 677.640 1747.000 679.640 ;
        RECT 4.400 676.240 1747.000 677.640 ;
        RECT 3.750 674.240 1747.000 676.240 ;
        RECT 4.400 672.840 1747.000 674.240 ;
        RECT 3.750 670.840 1747.000 672.840 ;
        RECT 4.400 669.440 1747.000 670.840 ;
        RECT 3.750 667.440 1747.000 669.440 ;
        RECT 4.400 666.040 1747.000 667.440 ;
        RECT 3.750 664.040 1747.000 666.040 ;
        RECT 4.400 662.640 1747.000 664.040 ;
        RECT 3.750 660.640 1747.000 662.640 ;
        RECT 4.400 659.240 1747.000 660.640 ;
        RECT 3.750 657.240 1747.000 659.240 ;
        RECT 4.400 655.840 1747.000 657.240 ;
        RECT 3.750 653.840 1747.000 655.840 ;
        RECT 4.400 652.440 1747.000 653.840 ;
        RECT 3.750 650.440 1747.000 652.440 ;
        RECT 4.400 649.040 1747.000 650.440 ;
        RECT 3.750 647.040 1747.000 649.040 ;
        RECT 4.400 645.640 1747.000 647.040 ;
        RECT 3.750 643.640 1747.000 645.640 ;
        RECT 4.400 642.240 1747.000 643.640 ;
        RECT 3.750 640.240 1747.000 642.240 ;
        RECT 4.400 638.840 1747.000 640.240 ;
        RECT 3.750 636.840 1747.000 638.840 ;
        RECT 4.400 635.440 1747.000 636.840 ;
        RECT 3.750 633.440 1747.000 635.440 ;
        RECT 4.400 632.040 1747.000 633.440 ;
        RECT 3.750 630.040 1747.000 632.040 ;
        RECT 4.400 628.640 1747.000 630.040 ;
        RECT 3.750 626.640 1747.000 628.640 ;
        RECT 4.400 625.240 1747.000 626.640 ;
        RECT 3.750 623.240 1747.000 625.240 ;
        RECT 4.400 621.840 1747.000 623.240 ;
        RECT 3.750 619.840 1747.000 621.840 ;
        RECT 4.400 618.440 1747.000 619.840 ;
        RECT 3.750 616.440 1747.000 618.440 ;
        RECT 4.400 615.040 1747.000 616.440 ;
        RECT 3.750 613.040 1747.000 615.040 ;
        RECT 4.400 611.640 1747.000 613.040 ;
        RECT 3.750 609.640 1747.000 611.640 ;
        RECT 4.400 608.240 1747.000 609.640 ;
        RECT 3.750 606.240 1747.000 608.240 ;
        RECT 4.400 604.840 1747.000 606.240 ;
        RECT 3.750 602.840 1747.000 604.840 ;
        RECT 4.400 601.440 1747.000 602.840 ;
        RECT 3.750 599.440 1747.000 601.440 ;
        RECT 4.400 598.040 1747.000 599.440 ;
        RECT 3.750 596.040 1747.000 598.040 ;
        RECT 4.400 594.640 1747.000 596.040 ;
        RECT 3.750 592.640 1747.000 594.640 ;
        RECT 4.400 591.240 1747.000 592.640 ;
        RECT 3.750 589.240 1747.000 591.240 ;
        RECT 4.400 587.840 1747.000 589.240 ;
        RECT 3.750 585.840 1747.000 587.840 ;
        RECT 4.400 584.440 1747.000 585.840 ;
        RECT 3.750 582.440 1747.000 584.440 ;
        RECT 4.400 581.040 1747.000 582.440 ;
        RECT 3.750 579.040 1747.000 581.040 ;
        RECT 4.400 577.640 1747.000 579.040 ;
        RECT 3.750 575.640 1747.000 577.640 ;
        RECT 4.400 574.240 1747.000 575.640 ;
        RECT 3.750 572.240 1747.000 574.240 ;
        RECT 4.400 570.840 1747.000 572.240 ;
        RECT 3.750 568.840 1747.000 570.840 ;
        RECT 4.400 567.440 1747.000 568.840 ;
        RECT 3.750 565.440 1747.000 567.440 ;
        RECT 4.400 564.040 1747.000 565.440 ;
        RECT 3.750 562.040 1747.000 564.040 ;
        RECT 4.400 560.640 1747.000 562.040 ;
        RECT 3.750 558.640 1747.000 560.640 ;
        RECT 4.400 557.240 1747.000 558.640 ;
        RECT 3.750 555.240 1747.000 557.240 ;
        RECT 4.400 553.840 1747.000 555.240 ;
        RECT 3.750 551.840 1747.000 553.840 ;
        RECT 4.400 550.440 1747.000 551.840 ;
        RECT 3.750 548.440 1747.000 550.440 ;
        RECT 4.400 547.040 1747.000 548.440 ;
        RECT 3.750 10.715 1747.000 547.040 ;
      LAYER met4 ;
        RECT 3.975 20.575 20.640 1732.465 ;
        RECT 23.040 20.575 23.940 1732.465 ;
        RECT 26.340 20.575 174.240 1732.465 ;
        RECT 176.640 20.575 177.540 1732.465 ;
        RECT 179.940 20.575 327.840 1732.465 ;
        RECT 330.240 20.575 331.140 1732.465 ;
        RECT 333.540 20.575 481.440 1732.465 ;
        RECT 483.840 20.575 484.740 1732.465 ;
        RECT 487.140 20.575 635.040 1732.465 ;
        RECT 637.440 20.575 638.340 1732.465 ;
        RECT 640.740 20.575 788.640 1732.465 ;
        RECT 791.040 20.575 791.940 1732.465 ;
        RECT 794.340 20.575 928.905 1732.465 ;
  END
END systolic_sorter
END LIBRARY

