module systolic_sorter (clk,
    load,
    rst,
    in_data_flat,
    out_data_flat);
 input clk;
 input load;
 input rst;
 input [255:0] in_data_flat;
 output [255:0] out_data_flat;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire \gen_left[0][0] ;
 wire \gen_left[0][10] ;
 wire \gen_left[0][11] ;
 wire \gen_left[0][12] ;
 wire \gen_left[0][13] ;
 wire \gen_left[0][14] ;
 wire \gen_left[0][15] ;
 wire \gen_left[0][16] ;
 wire \gen_left[0][17] ;
 wire \gen_left[0][18] ;
 wire \gen_left[0][19] ;
 wire \gen_left[0][1] ;
 wire \gen_left[0][20] ;
 wire \gen_left[0][21] ;
 wire \gen_left[0][22] ;
 wire \gen_left[0][23] ;
 wire \gen_left[0][24] ;
 wire \gen_left[0][25] ;
 wire \gen_left[0][26] ;
 wire \gen_left[0][27] ;
 wire \gen_left[0][28] ;
 wire \gen_left[0][29] ;
 wire \gen_left[0][2] ;
 wire \gen_left[0][30] ;
 wire \gen_left[0][31] ;
 wire \gen_left[0][3] ;
 wire \gen_left[0][4] ;
 wire \gen_left[0][5] ;
 wire \gen_left[0][6] ;
 wire \gen_left[0][7] ;
 wire \gen_left[0][8] ;
 wire \gen_left[0][9] ;
 wire \gen_left[1][0] ;
 wire \gen_left[1][10] ;
 wire \gen_left[1][11] ;
 wire \gen_left[1][12] ;
 wire \gen_left[1][13] ;
 wire \gen_left[1][14] ;
 wire \gen_left[1][15] ;
 wire \gen_left[1][16] ;
 wire \gen_left[1][17] ;
 wire \gen_left[1][18] ;
 wire \gen_left[1][19] ;
 wire \gen_left[1][1] ;
 wire \gen_left[1][20] ;
 wire \gen_left[1][21] ;
 wire \gen_left[1][22] ;
 wire \gen_left[1][23] ;
 wire \gen_left[1][24] ;
 wire \gen_left[1][25] ;
 wire \gen_left[1][26] ;
 wire \gen_left[1][27] ;
 wire \gen_left[1][28] ;
 wire \gen_left[1][29] ;
 wire \gen_left[1][2] ;
 wire \gen_left[1][30] ;
 wire \gen_left[1][31] ;
 wire \gen_left[1][3] ;
 wire \gen_left[1][4] ;
 wire \gen_left[1][5] ;
 wire \gen_left[1][6] ;
 wire \gen_left[1][7] ;
 wire \gen_left[1][8] ;
 wire \gen_left[1][9] ;
 wire \gen_left[2][0] ;
 wire \gen_left[2][10] ;
 wire \gen_left[2][11] ;
 wire \gen_left[2][12] ;
 wire \gen_left[2][13] ;
 wire \gen_left[2][14] ;
 wire \gen_left[2][15] ;
 wire \gen_left[2][16] ;
 wire \gen_left[2][17] ;
 wire \gen_left[2][18] ;
 wire \gen_left[2][19] ;
 wire \gen_left[2][1] ;
 wire \gen_left[2][20] ;
 wire \gen_left[2][21] ;
 wire \gen_left[2][22] ;
 wire \gen_left[2][23] ;
 wire \gen_left[2][24] ;
 wire \gen_left[2][25] ;
 wire \gen_left[2][26] ;
 wire \gen_left[2][27] ;
 wire \gen_left[2][28] ;
 wire \gen_left[2][29] ;
 wire \gen_left[2][2] ;
 wire \gen_left[2][30] ;
 wire \gen_left[2][31] ;
 wire \gen_left[2][3] ;
 wire \gen_left[2][4] ;
 wire \gen_left[2][5] ;
 wire \gen_left[2][6] ;
 wire \gen_left[2][7] ;
 wire \gen_left[2][8] ;
 wire \gen_left[2][9] ;
 wire \gen_left[3][0] ;
 wire \gen_left[3][10] ;
 wire \gen_left[3][11] ;
 wire \gen_left[3][12] ;
 wire \gen_left[3][13] ;
 wire \gen_left[3][14] ;
 wire \gen_left[3][15] ;
 wire \gen_left[3][16] ;
 wire \gen_left[3][17] ;
 wire \gen_left[3][18] ;
 wire \gen_left[3][19] ;
 wire \gen_left[3][1] ;
 wire \gen_left[3][20] ;
 wire \gen_left[3][21] ;
 wire \gen_left[3][22] ;
 wire \gen_left[3][23] ;
 wire \gen_left[3][24] ;
 wire \gen_left[3][25] ;
 wire \gen_left[3][26] ;
 wire \gen_left[3][27] ;
 wire \gen_left[3][28] ;
 wire \gen_left[3][29] ;
 wire \gen_left[3][2] ;
 wire \gen_left[3][30] ;
 wire \gen_left[3][31] ;
 wire \gen_left[3][3] ;
 wire \gen_left[3][4] ;
 wire \gen_left[3][5] ;
 wire \gen_left[3][6] ;
 wire \gen_left[3][7] ;
 wire \gen_left[3][8] ;
 wire \gen_left[3][9] ;
 wire \gen_left[4][0] ;
 wire \gen_left[4][10] ;
 wire \gen_left[4][11] ;
 wire \gen_left[4][12] ;
 wire \gen_left[4][13] ;
 wire \gen_left[4][14] ;
 wire \gen_left[4][15] ;
 wire \gen_left[4][16] ;
 wire \gen_left[4][17] ;
 wire \gen_left[4][18] ;
 wire \gen_left[4][19] ;
 wire \gen_left[4][1] ;
 wire \gen_left[4][20] ;
 wire \gen_left[4][21] ;
 wire \gen_left[4][22] ;
 wire \gen_left[4][23] ;
 wire \gen_left[4][24] ;
 wire \gen_left[4][25] ;
 wire \gen_left[4][26] ;
 wire \gen_left[4][27] ;
 wire \gen_left[4][28] ;
 wire \gen_left[4][29] ;
 wire \gen_left[4][2] ;
 wire \gen_left[4][30] ;
 wire \gen_left[4][31] ;
 wire \gen_left[4][3] ;
 wire \gen_left[4][4] ;
 wire \gen_left[4][5] ;
 wire \gen_left[4][6] ;
 wire \gen_left[4][7] ;
 wire \gen_left[4][8] ;
 wire \gen_left[4][9] ;
 wire \gen_left[5][0] ;
 wire \gen_left[5][10] ;
 wire \gen_left[5][11] ;
 wire \gen_left[5][12] ;
 wire \gen_left[5][13] ;
 wire \gen_left[5][14] ;
 wire \gen_left[5][15] ;
 wire \gen_left[5][16] ;
 wire \gen_left[5][17] ;
 wire \gen_left[5][18] ;
 wire \gen_left[5][19] ;
 wire \gen_left[5][1] ;
 wire \gen_left[5][20] ;
 wire \gen_left[5][21] ;
 wire \gen_left[5][22] ;
 wire \gen_left[5][23] ;
 wire \gen_left[5][24] ;
 wire \gen_left[5][25] ;
 wire \gen_left[5][26] ;
 wire \gen_left[5][27] ;
 wire \gen_left[5][28] ;
 wire \gen_left[5][29] ;
 wire \gen_left[5][2] ;
 wire \gen_left[5][30] ;
 wire \gen_left[5][31] ;
 wire \gen_left[5][3] ;
 wire \gen_left[5][4] ;
 wire \gen_left[5][5] ;
 wire \gen_left[5][6] ;
 wire \gen_left[5][7] ;
 wire \gen_left[5][8] ;
 wire \gen_left[5][9] ;
 wire \gen_left[6][0] ;
 wire \gen_left[6][10] ;
 wire \gen_left[6][11] ;
 wire \gen_left[6][12] ;
 wire \gen_left[6][13] ;
 wire \gen_left[6][14] ;
 wire \gen_left[6][15] ;
 wire \gen_left[6][16] ;
 wire \gen_left[6][17] ;
 wire \gen_left[6][18] ;
 wire \gen_left[6][19] ;
 wire \gen_left[6][1] ;
 wire \gen_left[6][20] ;
 wire \gen_left[6][21] ;
 wire \gen_left[6][22] ;
 wire \gen_left[6][23] ;
 wire \gen_left[6][24] ;
 wire \gen_left[6][25] ;
 wire \gen_left[6][26] ;
 wire \gen_left[6][27] ;
 wire \gen_left[6][28] ;
 wire \gen_left[6][29] ;
 wire \gen_left[6][2] ;
 wire \gen_left[6][30] ;
 wire \gen_left[6][31] ;
 wire \gen_left[6][3] ;
 wire \gen_left[6][4] ;
 wire \gen_left[6][5] ;
 wire \gen_left[6][6] ;
 wire \gen_left[6][7] ;
 wire \gen_left[6][8] ;
 wire \gen_left[6][9] ;
 wire \gen_pe[0].pe_inst.out_right[0] ;
 wire \gen_pe[0].pe_inst.out_right[10] ;
 wire \gen_pe[0].pe_inst.out_right[11] ;
 wire \gen_pe[0].pe_inst.out_right[12] ;
 wire \gen_pe[0].pe_inst.out_right[13] ;
 wire \gen_pe[0].pe_inst.out_right[14] ;
 wire \gen_pe[0].pe_inst.out_right[15] ;
 wire \gen_pe[0].pe_inst.out_right[16] ;
 wire \gen_pe[0].pe_inst.out_right[17] ;
 wire \gen_pe[0].pe_inst.out_right[18] ;
 wire \gen_pe[0].pe_inst.out_right[19] ;
 wire \gen_pe[0].pe_inst.out_right[1] ;
 wire \gen_pe[0].pe_inst.out_right[20] ;
 wire \gen_pe[0].pe_inst.out_right[21] ;
 wire \gen_pe[0].pe_inst.out_right[22] ;
 wire \gen_pe[0].pe_inst.out_right[23] ;
 wire \gen_pe[0].pe_inst.out_right[24] ;
 wire \gen_pe[0].pe_inst.out_right[25] ;
 wire \gen_pe[0].pe_inst.out_right[26] ;
 wire \gen_pe[0].pe_inst.out_right[27] ;
 wire \gen_pe[0].pe_inst.out_right[28] ;
 wire \gen_pe[0].pe_inst.out_right[29] ;
 wire \gen_pe[0].pe_inst.out_right[2] ;
 wire \gen_pe[0].pe_inst.out_right[30] ;
 wire \gen_pe[0].pe_inst.out_right[31] ;
 wire \gen_pe[0].pe_inst.out_right[3] ;
 wire \gen_pe[0].pe_inst.out_right[4] ;
 wire \gen_pe[0].pe_inst.out_right[5] ;
 wire \gen_pe[0].pe_inst.out_right[6] ;
 wire \gen_pe[0].pe_inst.out_right[7] ;
 wire \gen_pe[0].pe_inst.out_right[8] ;
 wire \gen_pe[0].pe_inst.out_right[9] ;
 wire \gen_pe[1].pe_inst.out_right[0] ;
 wire \gen_pe[1].pe_inst.out_right[10] ;
 wire \gen_pe[1].pe_inst.out_right[11] ;
 wire \gen_pe[1].pe_inst.out_right[12] ;
 wire \gen_pe[1].pe_inst.out_right[13] ;
 wire \gen_pe[1].pe_inst.out_right[14] ;
 wire \gen_pe[1].pe_inst.out_right[15] ;
 wire \gen_pe[1].pe_inst.out_right[16] ;
 wire \gen_pe[1].pe_inst.out_right[17] ;
 wire \gen_pe[1].pe_inst.out_right[18] ;
 wire \gen_pe[1].pe_inst.out_right[19] ;
 wire \gen_pe[1].pe_inst.out_right[1] ;
 wire \gen_pe[1].pe_inst.out_right[20] ;
 wire \gen_pe[1].pe_inst.out_right[21] ;
 wire \gen_pe[1].pe_inst.out_right[22] ;
 wire \gen_pe[1].pe_inst.out_right[23] ;
 wire \gen_pe[1].pe_inst.out_right[24] ;
 wire \gen_pe[1].pe_inst.out_right[25] ;
 wire \gen_pe[1].pe_inst.out_right[26] ;
 wire \gen_pe[1].pe_inst.out_right[27] ;
 wire \gen_pe[1].pe_inst.out_right[28] ;
 wire \gen_pe[1].pe_inst.out_right[29] ;
 wire \gen_pe[1].pe_inst.out_right[2] ;
 wire \gen_pe[1].pe_inst.out_right[30] ;
 wire \gen_pe[1].pe_inst.out_right[31] ;
 wire \gen_pe[1].pe_inst.out_right[3] ;
 wire \gen_pe[1].pe_inst.out_right[4] ;
 wire \gen_pe[1].pe_inst.out_right[5] ;
 wire \gen_pe[1].pe_inst.out_right[6] ;
 wire \gen_pe[1].pe_inst.out_right[7] ;
 wire \gen_pe[1].pe_inst.out_right[8] ;
 wire \gen_pe[1].pe_inst.out_right[9] ;
 wire \gen_pe[1].pe_inst.sel ;
 wire \gen_pe[2].pe_inst.out_right[0] ;
 wire \gen_pe[2].pe_inst.out_right[10] ;
 wire \gen_pe[2].pe_inst.out_right[11] ;
 wire \gen_pe[2].pe_inst.out_right[12] ;
 wire \gen_pe[2].pe_inst.out_right[13] ;
 wire \gen_pe[2].pe_inst.out_right[14] ;
 wire \gen_pe[2].pe_inst.out_right[15] ;
 wire \gen_pe[2].pe_inst.out_right[16] ;
 wire \gen_pe[2].pe_inst.out_right[17] ;
 wire \gen_pe[2].pe_inst.out_right[18] ;
 wire \gen_pe[2].pe_inst.out_right[19] ;
 wire \gen_pe[2].pe_inst.out_right[1] ;
 wire \gen_pe[2].pe_inst.out_right[20] ;
 wire \gen_pe[2].pe_inst.out_right[21] ;
 wire \gen_pe[2].pe_inst.out_right[22] ;
 wire \gen_pe[2].pe_inst.out_right[23] ;
 wire \gen_pe[2].pe_inst.out_right[24] ;
 wire \gen_pe[2].pe_inst.out_right[25] ;
 wire \gen_pe[2].pe_inst.out_right[26] ;
 wire \gen_pe[2].pe_inst.out_right[27] ;
 wire \gen_pe[2].pe_inst.out_right[28] ;
 wire \gen_pe[2].pe_inst.out_right[29] ;
 wire \gen_pe[2].pe_inst.out_right[2] ;
 wire \gen_pe[2].pe_inst.out_right[30] ;
 wire \gen_pe[2].pe_inst.out_right[31] ;
 wire \gen_pe[2].pe_inst.out_right[3] ;
 wire \gen_pe[2].pe_inst.out_right[4] ;
 wire \gen_pe[2].pe_inst.out_right[5] ;
 wire \gen_pe[2].pe_inst.out_right[6] ;
 wire \gen_pe[2].pe_inst.out_right[7] ;
 wire \gen_pe[2].pe_inst.out_right[8] ;
 wire \gen_pe[2].pe_inst.out_right[9] ;
 wire \gen_pe[3].pe_inst.out_right[0] ;
 wire \gen_pe[3].pe_inst.out_right[10] ;
 wire \gen_pe[3].pe_inst.out_right[11] ;
 wire \gen_pe[3].pe_inst.out_right[12] ;
 wire \gen_pe[3].pe_inst.out_right[13] ;
 wire \gen_pe[3].pe_inst.out_right[14] ;
 wire \gen_pe[3].pe_inst.out_right[15] ;
 wire \gen_pe[3].pe_inst.out_right[16] ;
 wire \gen_pe[3].pe_inst.out_right[17] ;
 wire \gen_pe[3].pe_inst.out_right[18] ;
 wire \gen_pe[3].pe_inst.out_right[19] ;
 wire \gen_pe[3].pe_inst.out_right[1] ;
 wire \gen_pe[3].pe_inst.out_right[20] ;
 wire \gen_pe[3].pe_inst.out_right[21] ;
 wire \gen_pe[3].pe_inst.out_right[22] ;
 wire \gen_pe[3].pe_inst.out_right[23] ;
 wire \gen_pe[3].pe_inst.out_right[24] ;
 wire \gen_pe[3].pe_inst.out_right[25] ;
 wire \gen_pe[3].pe_inst.out_right[26] ;
 wire \gen_pe[3].pe_inst.out_right[27] ;
 wire \gen_pe[3].pe_inst.out_right[28] ;
 wire \gen_pe[3].pe_inst.out_right[29] ;
 wire \gen_pe[3].pe_inst.out_right[2] ;
 wire \gen_pe[3].pe_inst.out_right[30] ;
 wire \gen_pe[3].pe_inst.out_right[31] ;
 wire \gen_pe[3].pe_inst.out_right[3] ;
 wire \gen_pe[3].pe_inst.out_right[4] ;
 wire \gen_pe[3].pe_inst.out_right[5] ;
 wire \gen_pe[3].pe_inst.out_right[6] ;
 wire \gen_pe[3].pe_inst.out_right[7] ;
 wire \gen_pe[3].pe_inst.out_right[8] ;
 wire \gen_pe[3].pe_inst.out_right[9] ;
 wire \gen_pe[4].pe_inst.out_right[0] ;
 wire \gen_pe[4].pe_inst.out_right[10] ;
 wire \gen_pe[4].pe_inst.out_right[11] ;
 wire \gen_pe[4].pe_inst.out_right[12] ;
 wire \gen_pe[4].pe_inst.out_right[13] ;
 wire \gen_pe[4].pe_inst.out_right[14] ;
 wire \gen_pe[4].pe_inst.out_right[15] ;
 wire \gen_pe[4].pe_inst.out_right[16] ;
 wire \gen_pe[4].pe_inst.out_right[17] ;
 wire \gen_pe[4].pe_inst.out_right[18] ;
 wire \gen_pe[4].pe_inst.out_right[19] ;
 wire \gen_pe[4].pe_inst.out_right[1] ;
 wire \gen_pe[4].pe_inst.out_right[20] ;
 wire \gen_pe[4].pe_inst.out_right[21] ;
 wire \gen_pe[4].pe_inst.out_right[22] ;
 wire \gen_pe[4].pe_inst.out_right[23] ;
 wire \gen_pe[4].pe_inst.out_right[24] ;
 wire \gen_pe[4].pe_inst.out_right[25] ;
 wire \gen_pe[4].pe_inst.out_right[26] ;
 wire \gen_pe[4].pe_inst.out_right[27] ;
 wire \gen_pe[4].pe_inst.out_right[28] ;
 wire \gen_pe[4].pe_inst.out_right[29] ;
 wire \gen_pe[4].pe_inst.out_right[2] ;
 wire \gen_pe[4].pe_inst.out_right[30] ;
 wire \gen_pe[4].pe_inst.out_right[31] ;
 wire \gen_pe[4].pe_inst.out_right[3] ;
 wire \gen_pe[4].pe_inst.out_right[4] ;
 wire \gen_pe[4].pe_inst.out_right[5] ;
 wire \gen_pe[4].pe_inst.out_right[6] ;
 wire \gen_pe[4].pe_inst.out_right[7] ;
 wire \gen_pe[4].pe_inst.out_right[8] ;
 wire \gen_pe[4].pe_inst.out_right[9] ;
 wire \gen_pe[5].pe_inst.out_right[0] ;
 wire \gen_pe[5].pe_inst.out_right[10] ;
 wire \gen_pe[5].pe_inst.out_right[11] ;
 wire \gen_pe[5].pe_inst.out_right[12] ;
 wire \gen_pe[5].pe_inst.out_right[13] ;
 wire \gen_pe[5].pe_inst.out_right[14] ;
 wire \gen_pe[5].pe_inst.out_right[15] ;
 wire \gen_pe[5].pe_inst.out_right[16] ;
 wire \gen_pe[5].pe_inst.out_right[17] ;
 wire \gen_pe[5].pe_inst.out_right[18] ;
 wire \gen_pe[5].pe_inst.out_right[19] ;
 wire \gen_pe[5].pe_inst.out_right[1] ;
 wire \gen_pe[5].pe_inst.out_right[20] ;
 wire \gen_pe[5].pe_inst.out_right[21] ;
 wire \gen_pe[5].pe_inst.out_right[22] ;
 wire \gen_pe[5].pe_inst.out_right[23] ;
 wire \gen_pe[5].pe_inst.out_right[24] ;
 wire \gen_pe[5].pe_inst.out_right[25] ;
 wire \gen_pe[5].pe_inst.out_right[26] ;
 wire \gen_pe[5].pe_inst.out_right[27] ;
 wire \gen_pe[5].pe_inst.out_right[28] ;
 wire \gen_pe[5].pe_inst.out_right[29] ;
 wire \gen_pe[5].pe_inst.out_right[2] ;
 wire \gen_pe[5].pe_inst.out_right[30] ;
 wire \gen_pe[5].pe_inst.out_right[31] ;
 wire \gen_pe[5].pe_inst.out_right[3] ;
 wire \gen_pe[5].pe_inst.out_right[4] ;
 wire \gen_pe[5].pe_inst.out_right[5] ;
 wire \gen_pe[5].pe_inst.out_right[6] ;
 wire \gen_pe[5].pe_inst.out_right[7] ;
 wire \gen_pe[5].pe_inst.out_right[8] ;
 wire \gen_pe[5].pe_inst.out_right[9] ;
 wire \gen_pe[6].pe_inst.out_right[0] ;
 wire \gen_pe[6].pe_inst.out_right[10] ;
 wire \gen_pe[6].pe_inst.out_right[11] ;
 wire \gen_pe[6].pe_inst.out_right[12] ;
 wire \gen_pe[6].pe_inst.out_right[13] ;
 wire \gen_pe[6].pe_inst.out_right[14] ;
 wire \gen_pe[6].pe_inst.out_right[15] ;
 wire \gen_pe[6].pe_inst.out_right[16] ;
 wire \gen_pe[6].pe_inst.out_right[17] ;
 wire \gen_pe[6].pe_inst.out_right[18] ;
 wire \gen_pe[6].pe_inst.out_right[19] ;
 wire \gen_pe[6].pe_inst.out_right[1] ;
 wire \gen_pe[6].pe_inst.out_right[20] ;
 wire \gen_pe[6].pe_inst.out_right[21] ;
 wire \gen_pe[6].pe_inst.out_right[22] ;
 wire \gen_pe[6].pe_inst.out_right[23] ;
 wire \gen_pe[6].pe_inst.out_right[24] ;
 wire \gen_pe[6].pe_inst.out_right[25] ;
 wire \gen_pe[6].pe_inst.out_right[26] ;
 wire \gen_pe[6].pe_inst.out_right[27] ;
 wire \gen_pe[6].pe_inst.out_right[28] ;
 wire \gen_pe[6].pe_inst.out_right[29] ;
 wire \gen_pe[6].pe_inst.out_right[2] ;
 wire \gen_pe[6].pe_inst.out_right[30] ;
 wire \gen_pe[6].pe_inst.out_right[31] ;
 wire \gen_pe[6].pe_inst.out_right[3] ;
 wire \gen_pe[6].pe_inst.out_right[4] ;
 wire \gen_pe[6].pe_inst.out_right[5] ;
 wire \gen_pe[6].pe_inst.out_right[6] ;
 wire \gen_pe[6].pe_inst.out_right[7] ;
 wire \gen_pe[6].pe_inst.out_right[8] ;
 wire \gen_pe[6].pe_inst.out_right[9] ;

 sky130_fd_sc_hd__mux2_1 _2371_ (.A0(out_data_flat[167]),
    .A1(out_data_flat[135]),
    .S(_2106_),
    .X(_0478_));
 sky130_fd_sc_hd__mux2_1 _2372_ (.A0(out_data_flat[168]),
    .A1(out_data_flat[136]),
    .S(_2106_),
    .X(_0479_));
 sky130_fd_sc_hd__mux2_1 _2373_ (.A0(out_data_flat[169]),
    .A1(out_data_flat[137]),
    .S(_2106_),
    .X(_0480_));
 sky130_fd_sc_hd__mux2_1 _2374_ (.A0(out_data_flat[170]),
    .A1(out_data_flat[138]),
    .S(_2106_),
    .X(_0450_));
 sky130_fd_sc_hd__mux2_1 _2375_ (.A0(out_data_flat[171]),
    .A1(out_data_flat[139]),
    .S(_2106_),
    .X(_0451_));
 sky130_fd_sc_hd__mux2_1 _2376_ (.A0(out_data_flat[172]),
    .A1(out_data_flat[140]),
    .S(_2106_),
    .X(_0452_));
 sky130_fd_sc_hd__mux2_1 _2377_ (.A0(out_data_flat[173]),
    .A1(out_data_flat[141]),
    .S(_2106_),
    .X(_0453_));
 sky130_fd_sc_hd__mux2_1 _2378_ (.A0(out_data_flat[174]),
    .A1(out_data_flat[142]),
    .S(_2106_),
    .X(_0454_));
 sky130_fd_sc_hd__mux2_1 _2379_ (.A0(out_data_flat[175]),
    .A1(out_data_flat[143]),
    .S(_2106_),
    .X(_0455_));
 sky130_fd_sc_hd__mux2_1 _2380_ (.A0(out_data_flat[176]),
    .A1(out_data_flat[144]),
    .S(_2106_),
    .X(_0456_));
 sky130_fd_sc_hd__mux2_1 _2381_ (.A0(out_data_flat[177]),
    .A1(out_data_flat[145]),
    .S(_2106_),
    .X(_0457_));
 sky130_fd_sc_hd__mux2_1 _2382_ (.A0(out_data_flat[178]),
    .A1(out_data_flat[146]),
    .S(_2106_),
    .X(_0458_));
 sky130_fd_sc_hd__mux2_1 _2383_ (.A0(out_data_flat[179]),
    .A1(out_data_flat[147]),
    .S(_2106_),
    .X(_0459_));
 sky130_fd_sc_hd__mux2_1 _2384_ (.A0(out_data_flat[180]),
    .A1(out_data_flat[148]),
    .S(_2106_),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_1 _2385_ (.A0(out_data_flat[181]),
    .A1(out_data_flat[149]),
    .S(_2106_),
    .X(_0462_));
 sky130_fd_sc_hd__mux2_1 _2386_ (.A0(out_data_flat[182]),
    .A1(out_data_flat[150]),
    .S(_2106_),
    .X(_0463_));
 sky130_fd_sc_hd__mux2_1 _2387_ (.A0(out_data_flat[183]),
    .A1(out_data_flat[151]),
    .S(_2106_),
    .X(_0464_));
 sky130_fd_sc_hd__mux2_1 _2388_ (.A0(out_data_flat[184]),
    .A1(out_data_flat[152]),
    .S(_2106_),
    .X(_0465_));
 sky130_fd_sc_hd__mux2_1 _2389_ (.A0(out_data_flat[185]),
    .A1(out_data_flat[153]),
    .S(_2106_),
    .X(_0466_));
 sky130_fd_sc_hd__mux2_1 _2390_ (.A0(out_data_flat[186]),
    .A1(out_data_flat[154]),
    .S(_2106_),
    .X(_0467_));
 sky130_fd_sc_hd__mux2_1 _2391_ (.A0(out_data_flat[187]),
    .A1(out_data_flat[155]),
    .S(_2106_),
    .X(_0468_));
 sky130_fd_sc_hd__mux2_1 _2392_ (.A0(out_data_flat[188]),
    .A1(out_data_flat[156]),
    .S(_2106_),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_1 _2393_ (.A0(out_data_flat[189]),
    .A1(out_data_flat[157]),
    .S(_2106_),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _2394_ (.A0(out_data_flat[190]),
    .A1(out_data_flat[158]),
    .S(_2106_),
    .X(_0472_));
 sky130_fd_sc_hd__o21a_2 _2395_ (.A1(\gen_pe[1].pe_inst.sel ),
    .A2(out_data_flat[191]),
    .B1(out_data_flat[159]),
    .X(_0473_));
 sky130_fd_sc_hd__mux2_1 _2396_ (.A0(out_data_flat[128]),
    .A1(out_data_flat[160]),
    .S(_2106_),
    .X(_0481_));
 sky130_fd_sc_hd__mux2_1 _2397_ (.A0(out_data_flat[129]),
    .A1(out_data_flat[161]),
    .S(_2106_),
    .X(_0492_));
 sky130_fd_sc_hd__mux2_1 _2398_ (.A0(out_data_flat[130]),
    .A1(out_data_flat[162]),
    .S(_2106_),
    .X(_0503_));
 sky130_fd_sc_hd__mux2_1 _2399_ (.A0(out_data_flat[131]),
    .A1(out_data_flat[163]),
    .S(_2106_),
    .X(_0506_));
 sky130_fd_sc_hd__mux2_1 _2400_ (.A0(out_data_flat[132]),
    .A1(out_data_flat[164]),
    .S(_2106_),
    .X(_0507_));
 sky130_fd_sc_hd__mux2_1 _2401_ (.A0(out_data_flat[133]),
    .A1(out_data_flat[165]),
    .S(_2106_),
    .X(_0508_));
 sky130_fd_sc_hd__mux2_1 _2402_ (.A0(out_data_flat[134]),
    .A1(out_data_flat[166]),
    .S(_2106_),
    .X(_0509_));
 sky130_fd_sc_hd__mux2_1 _2403_ (.A0(out_data_flat[135]),
    .A1(out_data_flat[167]),
    .S(_2106_),
    .X(_0510_));
 sky130_fd_sc_hd__mux2_1 _2404_ (.A0(out_data_flat[136]),
    .A1(out_data_flat[168]),
    .S(_2106_),
    .X(_0511_));
 sky130_fd_sc_hd__mux2_1 _2405_ (.A0(out_data_flat[137]),
    .A1(out_data_flat[169]),
    .S(_2106_),
    .X(_0512_));
 sky130_fd_sc_hd__mux2_1 _2406_ (.A0(out_data_flat[138]),
    .A1(out_data_flat[170]),
    .S(_2106_),
    .X(_0482_));
 sky130_fd_sc_hd__mux2_1 _2407_ (.A0(out_data_flat[139]),
    .A1(out_data_flat[171]),
    .S(_2106_),
    .X(_0483_));
 sky130_fd_sc_hd__mux2_1 _2408_ (.A0(out_data_flat[140]),
    .A1(out_data_flat[172]),
    .S(_2106_),
    .X(_0484_));
 sky130_fd_sc_hd__mux2_1 _2409_ (.A0(out_data_flat[141]),
    .A1(out_data_flat[173]),
    .S(_2106_),
    .X(_0485_));
 sky130_fd_sc_hd__mux2_1 _2410_ (.A0(out_data_flat[142]),
    .A1(out_data_flat[174]),
    .S(_2106_),
    .X(_0486_));
 sky130_fd_sc_hd__mux2_1 _2411_ (.A0(out_data_flat[143]),
    .A1(out_data_flat[175]),
    .S(_2106_),
    .X(_0487_));
 sky130_fd_sc_hd__mux2_1 _2412_ (.A0(out_data_flat[144]),
    .A1(out_data_flat[176]),
    .S(_2106_),
    .X(_0488_));
 sky130_fd_sc_hd__mux2_1 _2413_ (.A0(out_data_flat[145]),
    .A1(out_data_flat[177]),
    .S(_2106_),
    .X(_0489_));
 sky130_fd_sc_hd__mux2_1 _2414_ (.A0(out_data_flat[146]),
    .A1(out_data_flat[178]),
    .S(_2106_),
    .X(_0490_));
 sky130_fd_sc_hd__mux2_1 _2415_ (.A0(out_data_flat[147]),
    .A1(out_data_flat[179]),
    .S(_2106_),
    .X(_0491_));
 sky130_fd_sc_hd__mux2_1 _2416_ (.A0(out_data_flat[148]),
    .A1(out_data_flat[180]),
    .S(_2106_),
    .X(_0493_));
 sky130_fd_sc_hd__mux2_1 _2417_ (.A0(out_data_flat[149]),
    .A1(out_data_flat[181]),
    .S(_2106_),
    .X(_0494_));
 sky130_fd_sc_hd__mux2_1 _2418_ (.A0(out_data_flat[150]),
    .A1(out_data_flat[182]),
    .S(_2106_),
    .X(_0495_));
 sky130_fd_sc_hd__mux2_1 _2419_ (.A0(out_data_flat[151]),
    .A1(out_data_flat[183]),
    .S(_2106_),
    .X(_0496_));
 sky130_fd_sc_hd__mux2_1 _2420_ (.A0(out_data_flat[152]),
    .A1(out_data_flat[184]),
    .S(_2106_),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_1 _2421_ (.A0(out_data_flat[153]),
    .A1(out_data_flat[185]),
    .S(_2106_),
    .X(_0498_));
 sky130_fd_sc_hd__mux2_1 _2422_ (.A0(out_data_flat[154]),
    .A1(out_data_flat[186]),
    .S(_2106_),
    .X(_0499_));
 sky130_fd_sc_hd__mux2_1 _2423_ (.A0(out_data_flat[155]),
    .A1(out_data_flat[187]),
    .S(_2106_),
    .X(_0500_));
 sky130_fd_sc_hd__mux2_1 _2424_ (.A0(out_data_flat[156]),
    .A1(out_data_flat[188]),
    .S(_2106_),
    .X(_0501_));
 sky130_fd_sc_hd__mux2_1 _2425_ (.A0(out_data_flat[157]),
    .A1(out_data_flat[189]),
    .S(_2106_),
    .X(_0502_));
 sky130_fd_sc_hd__mux2_1 _2426_ (.A0(out_data_flat[158]),
    .A1(out_data_flat[190]),
    .S(_2106_),
    .X(_0504_));
 sky130_fd_sc_hd__a21o_2 _2427_ (.A1(_1428_),
    .A2(out_data_flat[159]),
    .B1(out_data_flat[191]),
    .X(_0505_));
 sky130_fd_sc_hd__a22o_2 _2428_ (.A1(_1486_),
    .A2(out_data_flat[159]),
    .B1(out_data_flat[158]),
    .B2(_1487_),
    .X(_2107_));
 sky130_fd_sc_hd__nand2b_2 _2429_ (.A_N(out_data_flat[159]),
    .B(out_data_flat[127]),
    .Y(_2108_));
 sky130_fd_sc_hd__o221a_2 _2430_ (.A1(_1487_),
    .A2(out_data_flat[158]),
    .B1(out_data_flat[157]),
    .B2(_1488_),
    .C1(_2108_),
    .X(_2109_));
 sky130_fd_sc_hd__and2b_2 _2431_ (.A_N(_2107_),
    .B(_2109_),
    .X(_2110_));
 sky130_fd_sc_hd__nand2b_2 _2432_ (.A_N(out_data_flat[155]),
    .B(out_data_flat[123]),
    .Y(_2111_));
 sky130_fd_sc_hd__xnor2_2 _2433_ (.A(out_data_flat[122]),
    .B(out_data_flat[154]),
    .Y(_2112_));
 sky130_fd_sc_hd__o211a_2 _2434_ (.A1(_1492_),
    .A2(out_data_flat[153]),
    .B1(_2111_),
    .C1(_2112_),
    .X(_2113_));
 sky130_fd_sc_hd__nand2_2 _2435_ (.A(out_data_flat[124]),
    .B(_1522_),
    .Y(_2114_));
 sky130_fd_sc_hd__o221a_2 _2436_ (.A1(out_data_flat[123]),
    .A2(_1523_),
    .B1(out_data_flat[152]),
    .B2(_1493_),
    .C1(_2114_),
    .X(_2115_));
 sky130_fd_sc_hd__a22o_2 _2437_ (.A1(_1488_),
    .A2(out_data_flat[157]),
    .B1(out_data_flat[156]),
    .B2(_1489_),
    .X(_2116_));
 sky130_fd_sc_hd__a22o_2 _2438_ (.A1(_1492_),
    .A2(out_data_flat[153]),
    .B1(out_data_flat[152]),
    .B2(_1493_),
    .X(_2117_));
 sky130_fd_sc_hd__nor2_2 _2439_ (.A(_2116_),
    .B(_2117_),
    .Y(_2118_));
 sky130_fd_sc_hd__and4_2 _2440_ (.A(_2110_),
    .B(_2113_),
    .C(_2115_),
    .D(_2118_),
    .X(_2119_));
 sky130_fd_sc_hd__a22o_2 _2441_ (.A1(_1498_),
    .A2(out_data_flat[147]),
    .B1(out_data_flat[146]),
    .B2(_1499_),
    .X(_2120_));
 sky130_fd_sc_hd__o22a_2 _2442_ (.A1(_1499_),
    .A2(out_data_flat[146]),
    .B1(out_data_flat[145]),
    .B2(_1500_),
    .X(_2121_));
 sky130_fd_sc_hd__a22o_2 _2443_ (.A1(_1500_),
    .A2(out_data_flat[145]),
    .B1(out_data_flat[144]),
    .B2(_1501_),
    .X(_2122_));
 sky130_fd_sc_hd__a21o_2 _2444_ (.A1(_2121_),
    .A2(_2122_),
    .B1(_2120_),
    .X(_2123_));
 sky130_fd_sc_hd__nand2b_2 _2445_ (.A_N(out_data_flat[118]),
    .B(out_data_flat[150]),
    .Y(_2124_));
 sky130_fd_sc_hd__nand2b_2 _2446_ (.A_N(out_data_flat[117]),
    .B(out_data_flat[149]),
    .Y(_2125_));
 sky130_fd_sc_hd__nand2b_2 _2447_ (.A_N(out_data_flat[116]),
    .B(out_data_flat[148]),
    .Y(_2126_));
 sky130_fd_sc_hd__o2111a_2 _2448_ (.A1(out_data_flat[119]),
    .A2(_1525_),
    .B1(_2124_),
    .C1(_2125_),
    .D1(_2126_),
    .X(_2127_));
 sky130_fd_sc_hd__o22a_2 _2449_ (.A1(_1495_),
    .A2(out_data_flat[150]),
    .B1(out_data_flat[149]),
    .B2(_1496_),
    .X(_2128_));
 sky130_fd_sc_hd__nand2_2 _2450_ (.A(out_data_flat[119]),
    .B(_1525_),
    .Y(_2129_));
 sky130_fd_sc_hd__or2_2 _2451_ (.A(_1498_),
    .B(out_data_flat[147]),
    .X(_2130_));
 sky130_fd_sc_hd__o2111a_2 _2452_ (.A1(_1497_),
    .A2(out_data_flat[148]),
    .B1(_2127_),
    .C1(_2128_),
    .D1(_2129_),
    .X(_2131_));
 sky130_fd_sc_hd__nand3_2 _2453_ (.A(_2123_),
    .B(_2130_),
    .C(_2131_),
    .Y(_2132_));
 sky130_fd_sc_hd__a221o_2 _2454_ (.A1(_1494_),
    .A2(out_data_flat[151]),
    .B1(out_data_flat[150]),
    .B2(_1495_),
    .C1(_2128_),
    .X(_2133_));
 sky130_fd_sc_hd__nand2_2 _2455_ (.A(_2129_),
    .B(_2133_),
    .Y(_2134_));
 sky130_fd_sc_hd__o21ai_2 _2456_ (.A1(_2127_),
    .A2(_2134_),
    .B1(_2132_),
    .Y(_2135_));
 sky130_fd_sc_hd__and2b_2 _2457_ (.A_N(out_data_flat[110]),
    .B(out_data_flat[142]),
    .X(_2136_));
 sky130_fd_sc_hd__a21o_2 _2458_ (.A1(_1502_),
    .A2(out_data_flat[143]),
    .B1(_2136_),
    .X(_2137_));
 sky130_fd_sc_hd__and2b_2 _2459_ (.A_N(out_data_flat[109]),
    .B(out_data_flat[141]),
    .X(_2138_));
 sky130_fd_sc_hd__and2b_2 _2460_ (.A_N(out_data_flat[108]),
    .B(out_data_flat[140]),
    .X(_2139_));
 sky130_fd_sc_hd__a2111o_2 _2461_ (.A1(_1502_),
    .A2(out_data_flat[143]),
    .B1(_2136_),
    .C1(_2138_),
    .D1(_2139_),
    .X(_2140_));
 sky130_fd_sc_hd__a22oi_2 _2462_ (.A1(out_data_flat[110]),
    .A2(_1529_),
    .B1(_1530_),
    .B2(out_data_flat[109]),
    .Y(_2141_));
 sky130_fd_sc_hd__and2_2 _2463_ (.A(out_data_flat[108]),
    .B(_1531_),
    .X(_2142_));
 sky130_fd_sc_hd__or2_2 _2464_ (.A(_1502_),
    .B(out_data_flat[143]),
    .X(_2143_));
 sky130_fd_sc_hd__or4bb_2 _2465_ (.A(_2140_),
    .B(_2142_),
    .C_N(_2143_),
    .D_N(_2141_),
    .X(_2144_));
 sky130_fd_sc_hd__o22a_2 _2466_ (.A1(out_data_flat[107]),
    .A2(_1532_),
    .B1(_1533_),
    .B2(out_data_flat[106]),
    .X(_2145_));
 sky130_fd_sc_hd__and2_2 _2467_ (.A(out_data_flat[107]),
    .B(_1532_),
    .X(_2146_));
 sky130_fd_sc_hd__a22o_2 _2468_ (.A1(out_data_flat[106]),
    .A2(_1533_),
    .B1(_1534_),
    .B2(out_data_flat[105]),
    .X(_2147_));
 sky130_fd_sc_hd__or4b_2 _2469_ (.A(_2144_),
    .B(_2146_),
    .C(_2147_),
    .D_N(_2145_),
    .X(_2148_));
 sky130_fd_sc_hd__o22a_2 _2470_ (.A1(out_data_flat[105]),
    .A2(_1534_),
    .B1(_1535_),
    .B2(out_data_flat[104]),
    .X(_2149_));
 sky130_fd_sc_hd__and2_2 _2471_ (.A(out_data_flat[104]),
    .B(_1535_),
    .X(_2150_));
 sky130_fd_sc_hd__and2_2 _2472_ (.A(out_data_flat[103]),
    .B(_1536_),
    .X(_2151_));
 sky130_fd_sc_hd__o22a_2 _2473_ (.A1(out_data_flat[103]),
    .A2(_1536_),
    .B1(_1537_),
    .B2(out_data_flat[102]),
    .X(_2152_));
 sky130_fd_sc_hd__o2bb2a_2 _2474_ (.A1_N(_1503_),
    .A2_N(out_data_flat[133]),
    .B1(_1538_),
    .B2(out_data_flat[100]),
    .X(_2153_));
 sky130_fd_sc_hd__and2_2 _2475_ (.A(out_data_flat[102]),
    .B(_1537_),
    .X(_2154_));
 sky130_fd_sc_hd__nor2_2 _2476_ (.A(_1503_),
    .B(out_data_flat[133]),
    .Y(_2155_));
 sky130_fd_sc_hd__o31a_2 _2477_ (.A1(_2153_),
    .A2(_2154_),
    .A3(_2155_),
    .B1(_2152_),
    .X(_2156_));
 sky130_fd_sc_hd__o211a_2 _2478_ (.A1(out_data_flat[97]),
    .A2(_1541_),
    .B1(_1542_),
    .C1(out_data_flat[96]),
    .X(_2157_));
 sky130_fd_sc_hd__a22o_2 _2479_ (.A1(out_data_flat[98]),
    .A2(_1540_),
    .B1(_1541_),
    .B2(out_data_flat[97]),
    .X(_2158_));
 sky130_fd_sc_hd__o22a_2 _2480_ (.A1(out_data_flat[99]),
    .A2(_1539_),
    .B1(_1540_),
    .B2(out_data_flat[98]),
    .X(_2159_));
 sky130_fd_sc_hd__o21a_2 _2481_ (.A1(_2157_),
    .A2(_2158_),
    .B1(_2159_),
    .X(_2160_));
 sky130_fd_sc_hd__a221o_2 _2482_ (.A1(out_data_flat[100]),
    .A2(_1538_),
    .B1(_1539_),
    .B2(out_data_flat[99]),
    .C1(_2155_),
    .X(_2161_));
 sky130_fd_sc_hd__or4bb_2 _2483_ (.A(_2151_),
    .B(_2154_),
    .C_N(_2153_),
    .D_N(_2152_),
    .X(_2162_));
 sky130_fd_sc_hd__o32a_2 _2484_ (.A1(_2160_),
    .A2(_2161_),
    .A3(_2162_),
    .B1(_2156_),
    .B2(_2151_),
    .X(_2163_));
 sky130_fd_sc_hd__o211ai_2 _2485_ (.A1(_2137_),
    .A2(_2141_),
    .B1(_2143_),
    .C1(_2140_),
    .Y(_2164_));
 sky130_fd_sc_hd__or4b_2 _2486_ (.A(_2148_),
    .B(_2150_),
    .C(_2163_),
    .D_N(_2149_),
    .X(_2165_));
 sky130_fd_sc_hd__o32a_2 _2487_ (.A1(_2144_),
    .A2(_2145_),
    .A3(_2146_),
    .B1(_2148_),
    .B2(_2149_),
    .X(_2166_));
 sky130_fd_sc_hd__o221a_2 _2488_ (.A1(out_data_flat[113]),
    .A2(_1527_),
    .B1(_1528_),
    .B2(out_data_flat[112]),
    .C1(_2121_),
    .X(_2167_));
 sky130_fd_sc_hd__a21oi_2 _2489_ (.A1(out_data_flat[112]),
    .A2(_1528_),
    .B1(_2120_),
    .Y(_2168_));
 sky130_fd_sc_hd__and4_2 _2490_ (.A(_2130_),
    .B(_2131_),
    .C(_2167_),
    .D(_2168_),
    .X(_2169_));
 sky130_fd_sc_hd__nand2_2 _2491_ (.A(_2119_),
    .B(_2135_),
    .Y(_2170_));
 sky130_fd_sc_hd__nand2_2 _2492_ (.A(_2119_),
    .B(_2169_),
    .Y(_2171_));
 sky130_fd_sc_hd__a31o_2 _2493_ (.A1(_2164_),
    .A2(_2165_),
    .A3(_2166_),
    .B1(_2171_),
    .X(_2172_));
 sky130_fd_sc_hd__and3_2 _2494_ (.A(_1491_),
    .B(out_data_flat[154]),
    .C(_2111_),
    .X(_2173_));
 sky130_fd_sc_hd__a22o_2 _2495_ (.A1(_1490_),
    .A2(out_data_flat[155]),
    .B1(_2113_),
    .B2(_2117_),
    .X(_2174_));
 sky130_fd_sc_hd__o21a_2 _2496_ (.A1(_2173_),
    .A2(_2174_),
    .B1(_2114_),
    .X(_2175_));
 sky130_fd_sc_hd__o21a_2 _2497_ (.A1(_2116_),
    .A2(_2175_),
    .B1(_2110_),
    .X(_2176_));
 sky130_fd_sc_hd__a21oi_2 _2498_ (.A1(_2107_),
    .A2(_2108_),
    .B1(_2176_),
    .Y(_2177_));
 sky130_fd_sc_hd__and4_2 _2499_ (.A(\gen_pe[1].pe_inst.sel ),
    .B(_2170_),
    .C(_2172_),
    .D(_2177_),
    .X(_2178_));
 sky130_fd_sc_hd__mux2_1 _2500_ (.A0(out_data_flat[96]),
    .A1(out_data_flat[128]),
    .S(_2178_),
    .X(_0385_));
 sky130_fd_sc_hd__mux2_1 _2501_ (.A0(out_data_flat[97]),
    .A1(out_data_flat[129]),
    .S(_2178_),
    .X(_0396_));
 sky130_fd_sc_hd__mux2_1 _2502_ (.A0(out_data_flat[98]),
    .A1(out_data_flat[130]),
    .S(_2178_),
    .X(_0407_));
 sky130_fd_sc_hd__mux2_1 _2503_ (.A0(out_data_flat[99]),
    .A1(out_data_flat[131]),
    .S(_2178_),
    .X(_0410_));
 sky130_fd_sc_hd__mux2_1 _2504_ (.A0(out_data_flat[100]),
    .A1(out_data_flat[132]),
    .S(_2178_),
    .X(_0411_));
 sky130_fd_sc_hd__mux2_1 _2505_ (.A0(out_data_flat[101]),
    .A1(out_data_flat[133]),
    .S(_2178_),
    .X(_0412_));
 sky130_fd_sc_hd__mux2_1 _2506_ (.A0(out_data_flat[102]),
    .A1(out_data_flat[134]),
    .S(_2178_),
    .X(_0413_));
 sky130_fd_sc_hd__mux2_1 _2507_ (.A0(out_data_flat[103]),
    .A1(out_data_flat[135]),
    .S(_2178_),
    .X(_0414_));
 sky130_fd_sc_hd__mux2_1 _2508_ (.A0(out_data_flat[104]),
    .A1(out_data_flat[136]),
    .S(_2178_),
    .X(_0415_));
 sky130_fd_sc_hd__mux2_1 _2509_ (.A0(out_data_flat[105]),
    .A1(out_data_flat[137]),
    .S(_2178_),
    .X(_0416_));
 sky130_fd_sc_hd__mux2_1 _2510_ (.A0(out_data_flat[106]),
    .A1(out_data_flat[138]),
    .S(_2178_),
    .X(_0386_));
 sky130_fd_sc_hd__mux2_1 _2511_ (.A0(out_data_flat[107]),
    .A1(out_data_flat[139]),
    .S(_2178_),
    .X(_0387_));
 sky130_fd_sc_hd__mux2_1 _2512_ (.A0(out_data_flat[108]),
    .A1(out_data_flat[140]),
    .S(_2178_),
    .X(_0388_));
 sky130_fd_sc_hd__mux2_1 _2513_ (.A0(out_data_flat[109]),
    .A1(out_data_flat[141]),
    .S(_2178_),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_1 _2514_ (.A0(out_data_flat[110]),
    .A1(out_data_flat[142]),
    .S(_2178_),
    .X(_0390_));
 sky130_fd_sc_hd__mux2_1 _2515_ (.A0(out_data_flat[111]),
    .A1(out_data_flat[143]),
    .S(_2178_),
    .X(_0391_));
 sky130_fd_sc_hd__mux2_1 _2516_ (.A0(out_data_flat[112]),
    .A1(out_data_flat[144]),
    .S(_2178_),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_1 _2517_ (.A0(out_data_flat[113]),
    .A1(out_data_flat[145]),
    .S(_2178_),
    .X(_0393_));
 sky130_fd_sc_hd__mux2_1 _2518_ (.A0(out_data_flat[114]),
    .A1(out_data_flat[146]),
    .S(_2178_),
    .X(_0394_));
 sky130_fd_sc_hd__mux2_1 _2519_ (.A0(out_data_flat[115]),
    .A1(out_data_flat[147]),
    .S(_2178_),
    .X(_0395_));
 sky130_fd_sc_hd__mux2_1 _2520_ (.A0(out_data_flat[116]),
    .A1(out_data_flat[148]),
    .S(_2178_),
    .X(_0397_));
 sky130_fd_sc_hd__mux2_1 _2521_ (.A0(out_data_flat[117]),
    .A1(out_data_flat[149]),
    .S(_2178_),
    .X(_0398_));
 sky130_fd_sc_hd__mux2_1 _2522_ (.A0(out_data_flat[118]),
    .A1(out_data_flat[150]),
    .S(_2178_),
    .X(_0399_));
 sky130_fd_sc_hd__mux2_1 _2523_ (.A0(out_data_flat[119]),
    .A1(out_data_flat[151]),
    .S(_2178_),
    .X(_0400_));
 sky130_fd_sc_hd__mux2_1 _2524_ (.A0(out_data_flat[120]),
    .A1(out_data_flat[152]),
    .S(_2178_),
    .X(_0401_));
 sky130_fd_sc_hd__mux2_1 _2525_ (.A0(out_data_flat[121]),
    .A1(out_data_flat[153]),
    .S(_2178_),
    .X(_0402_));
 sky130_fd_sc_hd__mux2_1 _2526_ (.A0(out_data_flat[122]),
    .A1(out_data_flat[154]),
    .S(_2178_),
    .X(_0403_));
 sky130_fd_sc_hd__mux2_1 _2527_ (.A0(out_data_flat[123]),
    .A1(out_data_flat[155]),
    .S(_2178_),
    .X(_0404_));
 sky130_fd_sc_hd__mux2_1 _2528_ (.A0(out_data_flat[124]),
    .A1(out_data_flat[156]),
    .S(_2178_),
    .X(_0405_));
 sky130_fd_sc_hd__mux2_1 _2529_ (.A0(out_data_flat[125]),
    .A1(out_data_flat[157]),
    .S(_2178_),
    .X(_0406_));
 sky130_fd_sc_hd__mux2_1 _2530_ (.A0(out_data_flat[126]),
    .A1(out_data_flat[158]),
    .S(_2178_),
    .X(_0408_));
 sky130_fd_sc_hd__a21oi_2 _2531_ (.A1(\gen_pe[1].pe_inst.sel ),
    .A2(_1521_),
    .B1(_1486_),
    .Y(_0409_));
 sky130_fd_sc_hd__mux2_1 _2532_ (.A0(out_data_flat[128]),
    .A1(out_data_flat[96]),
    .S(_2178_),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _2533_ (.A0(out_data_flat[129]),
    .A1(out_data_flat[97]),
    .S(_2178_),
    .X(_0428_));
 sky130_fd_sc_hd__mux2_1 _2534_ (.A0(out_data_flat[130]),
    .A1(out_data_flat[98]),
    .S(_2178_),
    .X(_0439_));
 sky130_fd_sc_hd__mux2_1 _2535_ (.A0(out_data_flat[131]),
    .A1(out_data_flat[99]),
    .S(_2178_),
    .X(_0442_));
 sky130_fd_sc_hd__mux2_1 _2536_ (.A0(out_data_flat[132]),
    .A1(out_data_flat[100]),
    .S(_2178_),
    .X(_0443_));
 sky130_fd_sc_hd__mux2_1 _2537_ (.A0(out_data_flat[133]),
    .A1(out_data_flat[101]),
    .S(_2178_),
    .X(_0444_));
 sky130_fd_sc_hd__mux2_1 _2538_ (.A0(out_data_flat[134]),
    .A1(out_data_flat[102]),
    .S(_2178_),
    .X(_0445_));
 sky130_fd_sc_hd__mux2_1 _2539_ (.A0(out_data_flat[135]),
    .A1(out_data_flat[103]),
    .S(_2178_),
    .X(_0446_));
 sky130_fd_sc_hd__mux2_1 _2540_ (.A0(out_data_flat[136]),
    .A1(out_data_flat[104]),
    .S(_2178_),
    .X(_0447_));
 sky130_fd_sc_hd__mux2_1 _2541_ (.A0(out_data_flat[137]),
    .A1(out_data_flat[105]),
    .S(_2178_),
    .X(_0448_));
 sky130_fd_sc_hd__mux2_1 _2542_ (.A0(out_data_flat[138]),
    .A1(out_data_flat[106]),
    .S(_2178_),
    .X(_0418_));
 sky130_fd_sc_hd__mux2_1 _2543_ (.A0(out_data_flat[139]),
    .A1(out_data_flat[107]),
    .S(_2178_),
    .X(_0419_));
 sky130_fd_sc_hd__mux2_1 _2544_ (.A0(out_data_flat[140]),
    .A1(out_data_flat[108]),
    .S(_2178_),
    .X(_0420_));
 sky130_fd_sc_hd__mux2_1 _2545_ (.A0(out_data_flat[141]),
    .A1(out_data_flat[109]),
    .S(_2178_),
    .X(_0421_));
 sky130_fd_sc_hd__mux2_1 _2546_ (.A0(out_data_flat[142]),
    .A1(out_data_flat[110]),
    .S(_2178_),
    .X(_0422_));
 sky130_fd_sc_hd__mux2_1 _2547_ (.A0(out_data_flat[143]),
    .A1(out_data_flat[111]),
    .S(_2178_),
    .X(_0423_));
 sky130_fd_sc_hd__mux2_1 _2548_ (.A0(out_data_flat[144]),
    .A1(out_data_flat[112]),
    .S(_2178_),
    .X(_0424_));
 sky130_fd_sc_hd__mux2_1 _2549_ (.A0(out_data_flat[145]),
    .A1(out_data_flat[113]),
    .S(_2178_),
    .X(_0425_));
 sky130_fd_sc_hd__mux2_1 _2550_ (.A0(out_data_flat[146]),
    .A1(out_data_flat[114]),
    .S(_2178_),
    .X(_0426_));
 sky130_fd_sc_hd__mux2_1 _2551_ (.A0(out_data_flat[147]),
    .A1(out_data_flat[115]),
    .S(_2178_),
    .X(_0427_));
 sky130_fd_sc_hd__mux2_1 _2552_ (.A0(out_data_flat[148]),
    .A1(out_data_flat[116]),
    .S(_2178_),
    .X(_0429_));
 sky130_fd_sc_hd__mux2_1 _2553_ (.A0(out_data_flat[149]),
    .A1(out_data_flat[117]),
    .S(_2178_),
    .X(_0430_));
 sky130_fd_sc_hd__mux2_1 _2554_ (.A0(out_data_flat[150]),
    .A1(out_data_flat[118]),
    .S(_2178_),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_1 _2555_ (.A0(out_data_flat[151]),
    .A1(out_data_flat[119]),
    .S(_2178_),
    .X(_0432_));
 sky130_fd_sc_hd__mux2_1 _2556_ (.A0(out_data_flat[152]),
    .A1(out_data_flat[120]),
    .S(_2178_),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_1 _2557_ (.A0(out_data_flat[153]),
    .A1(out_data_flat[121]),
    .S(_2178_),
    .X(_0434_));
 sky130_fd_sc_hd__mux2_1 _2558_ (.A0(out_data_flat[154]),
    .A1(out_data_flat[122]),
    .S(_2178_),
    .X(_0435_));
 sky130_fd_sc_hd__mux2_1 _2559_ (.A0(out_data_flat[155]),
    .A1(out_data_flat[123]),
    .S(_2178_),
    .X(_0436_));
 sky130_fd_sc_hd__mux2_1 _2560_ (.A0(out_data_flat[156]),
    .A1(out_data_flat[124]),
    .S(_2178_),
    .X(_0437_));
 sky130_fd_sc_hd__mux2_1 _2561_ (.A0(out_data_flat[157]),
    .A1(out_data_flat[125]),
    .S(_2178_),
    .X(_0438_));
 sky130_fd_sc_hd__mux2_1 _2562_ (.A0(out_data_flat[158]),
    .A1(out_data_flat[126]),
    .S(_2178_),
    .X(_0440_));
 sky130_fd_sc_hd__a21o_2 _2563_ (.A1(\gen_pe[1].pe_inst.sel ),
    .A2(out_data_flat[127]),
    .B1(out_data_flat[159]),
    .X(_0441_));
 sky130_fd_sc_hd__mux2_1 _2564_ (.A0(out_data_flat[192]),
    .A1(out_data_flat[224]),
    .S(_1775_),
    .X(_0609_));
 sky130_fd_sc_hd__mux2_1 _2565_ (.A0(out_data_flat[193]),
    .A1(out_data_flat[225]),
    .S(_1775_),
    .X(_0620_));
 sky130_fd_sc_hd__mux2_1 _2566_ (.A0(out_data_flat[194]),
    .A1(out_data_flat[226]),
    .S(_1775_),
    .X(_0631_));
 sky130_fd_sc_hd__mux2_1 _2567_ (.A0(out_data_flat[195]),
    .A1(out_data_flat[227]),
    .S(_1775_),
    .X(_0634_));
 sky130_fd_sc_hd__mux2_1 _2568_ (.A0(out_data_flat[196]),
    .A1(out_data_flat[228]),
    .S(_1775_),
    .X(_0635_));
 sky130_fd_sc_hd__mux2_1 _2569_ (.A0(out_data_flat[197]),
    .A1(out_data_flat[229]),
    .S(_1775_),
    .X(_0636_));
 sky130_fd_sc_hd__mux2_1 _2570_ (.A0(out_data_flat[198]),
    .A1(out_data_flat[230]),
    .S(_1775_),
    .X(_0637_));
 sky130_fd_sc_hd__mux2_1 _2571_ (.A0(out_data_flat[199]),
    .A1(out_data_flat[231]),
    .S(_1775_),
    .X(_0638_));
 sky130_fd_sc_hd__mux2_1 _2572_ (.A0(out_data_flat[200]),
    .A1(out_data_flat[232]),
    .S(_1775_),
    .X(_0639_));
 sky130_fd_sc_hd__mux2_1 _2573_ (.A0(out_data_flat[201]),
    .A1(out_data_flat[233]),
    .S(_1775_),
    .X(_0640_));
 sky130_fd_sc_hd__mux2_1 _2574_ (.A0(out_data_flat[202]),
    .A1(out_data_flat[234]),
    .S(_1775_),
    .X(_0610_));
 sky130_fd_sc_hd__mux2_1 _2575_ (.A0(out_data_flat[203]),
    .A1(out_data_flat[235]),
    .S(_1775_),
    .X(_0611_));
 sky130_fd_sc_hd__mux2_1 _2576_ (.A0(out_data_flat[204]),
    .A1(out_data_flat[236]),
    .S(_1775_),
    .X(_0612_));
 sky130_fd_sc_hd__mux2_1 _2577_ (.A0(out_data_flat[205]),
    .A1(out_data_flat[237]),
    .S(_1775_),
    .X(_0613_));
 sky130_fd_sc_hd__mux2_1 _2578_ (.A0(out_data_flat[206]),
    .A1(out_data_flat[238]),
    .S(_1775_),
    .X(_0614_));
 sky130_fd_sc_hd__mux2_1 _2579_ (.A0(out_data_flat[207]),
    .A1(out_data_flat[239]),
    .S(_1775_),
    .X(_0615_));
 sky130_fd_sc_hd__mux2_1 _2580_ (.A0(out_data_flat[208]),
    .A1(out_data_flat[240]),
    .S(_1775_),
    .X(_0616_));
 sky130_fd_sc_hd__mux2_1 _2581_ (.A0(out_data_flat[209]),
    .A1(out_data_flat[241]),
    .S(_1775_),
    .X(_0617_));
 sky130_fd_sc_hd__mux2_1 _2582_ (.A0(out_data_flat[210]),
    .A1(out_data_flat[242]),
    .S(_1775_),
    .X(_0618_));
 sky130_fd_sc_hd__mux2_1 _2583_ (.A0(out_data_flat[211]),
    .A1(out_data_flat[243]),
    .S(_1775_),
    .X(_0619_));
 sky130_fd_sc_hd__mux2_1 _2584_ (.A0(out_data_flat[212]),
    .A1(out_data_flat[244]),
    .S(_1775_),
    .X(_0621_));
 sky130_fd_sc_hd__mux2_1 _2585_ (.A0(out_data_flat[213]),
    .A1(out_data_flat[245]),
    .S(_1775_),
    .X(_0622_));
 sky130_fd_sc_hd__mux2_1 _2586_ (.A0(out_data_flat[214]),
    .A1(out_data_flat[246]),
    .S(_1775_),
    .X(_0623_));
 sky130_fd_sc_hd__mux2_1 _2587_ (.A0(out_data_flat[215]),
    .A1(out_data_flat[247]),
    .S(_1775_),
    .X(_0624_));
 sky130_fd_sc_hd__mux2_1 _2588_ (.A0(out_data_flat[216]),
    .A1(out_data_flat[248]),
    .S(_1775_),
    .X(_0625_));
 sky130_fd_sc_hd__mux2_1 _2589_ (.A0(out_data_flat[217]),
    .A1(out_data_flat[249]),
    .S(_1775_),
    .X(_0626_));
 sky130_fd_sc_hd__mux2_1 _2590_ (.A0(out_data_flat[218]),
    .A1(out_data_flat[250]),
    .S(_1775_),
    .X(_0627_));
 sky130_fd_sc_hd__mux2_1 _2591_ (.A0(out_data_flat[219]),
    .A1(out_data_flat[251]),
    .S(_1775_),
    .X(_0628_));
 sky130_fd_sc_hd__mux2_1 _2592_ (.A0(out_data_flat[220]),
    .A1(out_data_flat[252]),
    .S(_1775_),
    .X(_0629_));
 sky130_fd_sc_hd__mux2_1 _2593_ (.A0(out_data_flat[221]),
    .A1(out_data_flat[253]),
    .S(_1775_),
    .X(_0630_));
 sky130_fd_sc_hd__mux2_1 _2594_ (.A0(out_data_flat[222]),
    .A1(out_data_flat[254]),
    .S(_1775_),
    .X(_0632_));
 sky130_fd_sc_hd__a21o_2 _2595_ (.A1(_1428_),
    .A2(out_data_flat[223]),
    .B1(out_data_flat[255]),
    .X(_0633_));
 sky130_fd_sc_hd__a22o_2 _2596_ (.A1(load),
    .A2(in_data_flat[32]),
    .B1(_0192_),
    .B2(\gen_pe[0].pe_inst.out_right[0] ),
    .X(_2179_));
 sky130_fd_sc_hd__a21o_2 _2597_ (.A1(\gen_left[1][0] ),
    .A2(_1543_),
    .B1(_2179_),
    .X(_0000_));
 sky130_fd_sc_hd__a22o_2 _2598_ (.A1(load),
    .A2(in_data_flat[33]),
    .B1(_0192_),
    .B2(\gen_pe[0].pe_inst.out_right[1] ),
    .X(_2180_));
 sky130_fd_sc_hd__a21o_2 _2599_ (.A1(\gen_left[1][1] ),
    .A2(_1543_),
    .B1(_2180_),
    .X(_0011_));
 sky130_fd_sc_hd__a22o_2 _2600_ (.A1(load),
    .A2(in_data_flat[34]),
    .B1(_0192_),
    .B2(\gen_pe[0].pe_inst.out_right[2] ),
    .X(_2181_));
 sky130_fd_sc_hd__a21o_2 _2601_ (.A1(\gen_left[1][2] ),
    .A2(_1543_),
    .B1(_2181_),
    .X(_0022_));
 sky130_fd_sc_hd__a22o_2 _2602_ (.A1(load),
    .A2(in_data_flat[35]),
    .B1(_0192_),
    .B2(\gen_pe[0].pe_inst.out_right[3] ),
    .X(_2182_));
 sky130_fd_sc_hd__a21o_2 _2603_ (.A1(\gen_left[1][3] ),
    .A2(_1543_),
    .B1(_2182_),
    .X(_0025_));
 sky130_fd_sc_hd__a22o_2 _2604_ (.A1(load),
    .A2(in_data_flat[36]),
    .B1(_0192_),
    .B2(\gen_pe[0].pe_inst.out_right[4] ),
    .X(_2183_));
 sky130_fd_sc_hd__a21o_2 _2605_ (.A1(\gen_left[1][4] ),
    .A2(_1543_),
    .B1(_2183_),
    .X(_0026_));
 sky130_fd_sc_hd__a22o_2 _2606_ (.A1(load),
    .A2(in_data_flat[37]),
    .B1(_0192_),
    .B2(\gen_pe[0].pe_inst.out_right[5] ),
    .X(_2184_));
 sky130_fd_sc_hd__a21o_2 _2607_ (.A1(\gen_left[1][5] ),
    .A2(_1543_),
    .B1(_2184_),
    .X(_0027_));
 sky130_fd_sc_hd__a22o_2 _2608_ (.A1(load),
    .A2(in_data_flat[38]),
    .B1(_0192_),
    .B2(\gen_pe[0].pe_inst.out_right[6] ),
    .X(_2185_));
 sky130_fd_sc_hd__a21o_2 _2609_ (.A1(\gen_left[1][6] ),
    .A2(_1543_),
    .B1(_2185_),
    .X(_0028_));
 sky130_fd_sc_hd__and2_2 _2610_ (.A(load),
    .B(in_data_flat[39]),
    .X(_2186_));
 sky130_fd_sc_hd__a221o_2 _2611_ (.A1(\gen_pe[0].pe_inst.out_right[7] ),
    .A2(_0192_),
    .B1(_1543_),
    .B2(\gen_left[1][7] ),
    .C1(_2186_),
    .X(_0029_));
 sky130_fd_sc_hd__a22o_2 _2612_ (.A1(load),
    .A2(in_data_flat[40]),
    .B1(_0192_),
    .B2(\gen_pe[0].pe_inst.out_right[8] ),
    .X(_2187_));
 sky130_fd_sc_hd__a21o_2 _2613_ (.A1(\gen_left[1][8] ),
    .A2(_1543_),
    .B1(_2187_),
    .X(_0030_));
 sky130_fd_sc_hd__a22o_2 _2614_ (.A1(load),
    .A2(in_data_flat[41]),
    .B1(_0192_),
    .B2(\gen_pe[0].pe_inst.out_right[9] ),
    .X(_2188_));
 sky130_fd_sc_hd__a21o_2 _2615_ (.A1(\gen_left[1][9] ),
    .A2(_1543_),
    .B1(_2188_),
    .X(_0031_));
 sky130_fd_sc_hd__a22o_2 _2616_ (.A1(load),
    .A2(in_data_flat[42]),
    .B1(_0192_),
    .B2(\gen_pe[0].pe_inst.out_right[10] ),
    .X(_2189_));
 sky130_fd_sc_hd__a21o_2 _2617_ (.A1(\gen_left[1][10] ),
    .A2(_1543_),
    .B1(_2189_),
    .X(_0001_));
 sky130_fd_sc_hd__a22o_2 _2618_ (.A1(load),
    .A2(in_data_flat[43]),
    .B1(_0192_),
    .B2(\gen_pe[0].pe_inst.out_right[11] ),
    .X(_2190_));
 sky130_fd_sc_hd__a21o_2 _2619_ (.A1(\gen_left[1][11] ),
    .A2(_1543_),
    .B1(_2190_),
    .X(_0002_));
 sky130_fd_sc_hd__a22o_2 _2620_ (.A1(load),
    .A2(in_data_flat[44]),
    .B1(_0192_),
    .B2(\gen_pe[0].pe_inst.out_right[12] ),
    .X(_2191_));
 sky130_fd_sc_hd__a21o_2 _2621_ (.A1(\gen_left[1][12] ),
    .A2(_1543_),
    .B1(_2191_),
    .X(_0003_));
 sky130_fd_sc_hd__a22o_2 _2622_ (.A1(load),
    .A2(in_data_flat[45]),
    .B1(_0192_),
    .B2(\gen_pe[0].pe_inst.out_right[13] ),
    .X(_2192_));
 sky130_fd_sc_hd__a21o_2 _2623_ (.A1(\gen_left[1][13] ),
    .A2(_1543_),
    .B1(_2192_),
    .X(_0004_));
 sky130_fd_sc_hd__and2_2 _2624_ (.A(load),
    .B(in_data_flat[46]),
    .X(_2193_));
 sky130_fd_sc_hd__a221o_2 _2625_ (.A1(\gen_pe[0].pe_inst.out_right[14] ),
    .A2(_0192_),
    .B1(_1543_),
    .B2(\gen_left[1][14] ),
    .C1(_2193_),
    .X(_0005_));
 sky130_fd_sc_hd__and2_2 _2626_ (.A(load),
    .B(in_data_flat[47]),
    .X(_2194_));
 sky130_fd_sc_hd__a221o_2 _2627_ (.A1(\gen_pe[0].pe_inst.out_right[15] ),
    .A2(_0192_),
    .B1(_1543_),
    .B2(\gen_left[1][15] ),
    .C1(_2194_),
    .X(_0006_));
 sky130_fd_sc_hd__a22o_2 _2628_ (.A1(load),
    .A2(in_data_flat[48]),
    .B1(_0192_),
    .B2(\gen_pe[0].pe_inst.out_right[16] ),
    .X(_2195_));
 sky130_fd_sc_hd__a21o_2 _2629_ (.A1(\gen_left[1][16] ),
    .A2(_1543_),
    .B1(_2195_),
    .X(_0007_));
 sky130_fd_sc_hd__a22o_2 _2630_ (.A1(load),
    .A2(in_data_flat[49]),
    .B1(_0192_),
    .B2(\gen_pe[0].pe_inst.out_right[17] ),
    .X(_2196_));
 sky130_fd_sc_hd__a21o_2 _2631_ (.A1(\gen_left[1][17] ),
    .A2(_1543_),
    .B1(_2196_),
    .X(_0008_));
 sky130_fd_sc_hd__a22o_2 _2632_ (.A1(load),
    .A2(in_data_flat[50]),
    .B1(_0192_),
    .B2(\gen_pe[0].pe_inst.out_right[18] ),
    .X(_2197_));
 sky130_fd_sc_hd__a21o_2 _2633_ (.A1(\gen_left[1][18] ),
    .A2(_1543_),
    .B1(_2197_),
    .X(_0009_));
 sky130_fd_sc_hd__a22o_2 _2634_ (.A1(load),
    .A2(in_data_flat[51]),
    .B1(_0192_),
    .B2(\gen_pe[0].pe_inst.out_right[19] ),
    .X(_2198_));
 sky130_fd_sc_hd__a21o_2 _2635_ (.A1(\gen_left[1][19] ),
    .A2(_1543_),
    .B1(_2198_),
    .X(_0010_));
 sky130_fd_sc_hd__a22o_2 _2636_ (.A1(load),
    .A2(in_data_flat[52]),
    .B1(_0192_),
    .B2(\gen_pe[0].pe_inst.out_right[20] ),
    .X(_2199_));
 sky130_fd_sc_hd__a21o_2 _2637_ (.A1(\gen_left[1][20] ),
    .A2(_1543_),
    .B1(_2199_),
    .X(_0012_));
 sky130_fd_sc_hd__a22o_2 _2638_ (.A1(load),
    .A2(in_data_flat[53]),
    .B1(_0192_),
    .B2(\gen_pe[0].pe_inst.out_right[21] ),
    .X(_2200_));
 sky130_fd_sc_hd__a21o_2 _2639_ (.A1(\gen_left[1][21] ),
    .A2(_1543_),
    .B1(_2200_),
    .X(_0013_));
 sky130_fd_sc_hd__a22o_2 _2640_ (.A1(load),
    .A2(in_data_flat[54]),
    .B1(_0192_),
    .B2(\gen_pe[0].pe_inst.out_right[22] ),
    .X(_2201_));
 sky130_fd_sc_hd__a21o_2 _2641_ (.A1(\gen_left[1][22] ),
    .A2(_1543_),
    .B1(_2201_),
    .X(_0014_));
 sky130_fd_sc_hd__a22o_2 _2642_ (.A1(load),
    .A2(in_data_flat[55]),
    .B1(_0192_),
    .B2(\gen_pe[0].pe_inst.out_right[23] ),
    .X(_2202_));
 sky130_fd_sc_hd__a21o_2 _2643_ (.A1(\gen_left[1][23] ),
    .A2(_1543_),
    .B1(_2202_),
    .X(_0015_));
 sky130_fd_sc_hd__a22o_2 _2644_ (.A1(load),
    .A2(in_data_flat[56]),
    .B1(_0192_),
    .B2(\gen_pe[0].pe_inst.out_right[24] ),
    .X(_2203_));
 sky130_fd_sc_hd__a21o_2 _2645_ (.A1(\gen_left[1][24] ),
    .A2(_1543_),
    .B1(_2203_),
    .X(_0016_));
 sky130_fd_sc_hd__and2_2 _2646_ (.A(load),
    .B(in_data_flat[57]),
    .X(_2204_));
 sky130_fd_sc_hd__a221o_2 _2647_ (.A1(\gen_pe[0].pe_inst.out_right[25] ),
    .A2(_0192_),
    .B1(_1543_),
    .B2(\gen_left[1][25] ),
    .C1(_2204_),
    .X(_0017_));
 sky130_fd_sc_hd__a22o_2 _2648_ (.A1(load),
    .A2(in_data_flat[58]),
    .B1(_0192_),
    .B2(\gen_pe[0].pe_inst.out_right[26] ),
    .X(_2205_));
 sky130_fd_sc_hd__a21o_2 _2649_ (.A1(\gen_left[1][26] ),
    .A2(_1543_),
    .B1(_2205_),
    .X(_0018_));
 sky130_fd_sc_hd__a22o_2 _2650_ (.A1(load),
    .A2(in_data_flat[59]),
    .B1(_0192_),
    .B2(\gen_pe[0].pe_inst.out_right[27] ),
    .X(_2206_));
 sky130_fd_sc_hd__a21o_2 _2651_ (.A1(\gen_left[1][27] ),
    .A2(_1543_),
    .B1(_2206_),
    .X(_0019_));
 sky130_fd_sc_hd__and2_2 _2652_ (.A(load),
    .B(in_data_flat[60]),
    .X(_2207_));
 sky130_fd_sc_hd__a221o_2 _2653_ (.A1(\gen_pe[0].pe_inst.out_right[28] ),
    .A2(_0192_),
    .B1(_1543_),
    .B2(\gen_left[1][28] ),
    .C1(_2207_),
    .X(_0020_));
 sky130_fd_sc_hd__a22o_2 _2654_ (.A1(load),
    .A2(in_data_flat[61]),
    .B1(_0192_),
    .B2(\gen_pe[0].pe_inst.out_right[29] ),
    .X(_2208_));
 sky130_fd_sc_hd__a21o_2 _2655_ (.A1(\gen_left[1][29] ),
    .A2(_1543_),
    .B1(_2208_),
    .X(_0021_));
 sky130_fd_sc_hd__a22o_2 _2656_ (.A1(load),
    .A2(in_data_flat[62]),
    .B1(_0192_),
    .B2(\gen_pe[0].pe_inst.out_right[30] ),
    .X(_2209_));
 sky130_fd_sc_hd__a21o_2 _2657_ (.A1(\gen_left[1][30] ),
    .A2(_1543_),
    .B1(_2209_),
    .X(_0023_));
 sky130_fd_sc_hd__a22o_2 _2658_ (.A1(load),
    .A2(in_data_flat[63]),
    .B1(_0192_),
    .B2(\gen_pe[0].pe_inst.out_right[31] ),
    .X(_2210_));
 sky130_fd_sc_hd__a21o_2 _2659_ (.A1(\gen_left[1][31] ),
    .A2(_1543_),
    .B1(_2210_),
    .X(_0024_));
 sky130_fd_sc_hd__a22o_2 _2660_ (.A1(load),
    .A2(in_data_flat[64]),
    .B1(_0192_),
    .B2(\gen_left[2][0] ),
    .X(_2211_));
 sky130_fd_sc_hd__a21o_2 _2661_ (.A1(\gen_pe[1].pe_inst.out_right[0] ),
    .A2(_1543_),
    .B1(_2211_),
    .X(_0032_));
 sky130_fd_sc_hd__a22o_2 _2662_ (.A1(load),
    .A2(in_data_flat[65]),
    .B1(_0192_),
    .B2(\gen_left[2][1] ),
    .X(_2212_));
 sky130_fd_sc_hd__a21o_2 _2663_ (.A1(\gen_pe[1].pe_inst.out_right[1] ),
    .A2(_1543_),
    .B1(_2212_),
    .X(_0043_));
 sky130_fd_sc_hd__a22o_2 _2664_ (.A1(load),
    .A2(in_data_flat[66]),
    .B1(_0192_),
    .B2(\gen_left[2][2] ),
    .X(_2213_));
 sky130_fd_sc_hd__a21o_2 _2665_ (.A1(\gen_pe[1].pe_inst.out_right[2] ),
    .A2(_1543_),
    .B1(_2213_),
    .X(_0054_));
 sky130_fd_sc_hd__a22o_2 _2666_ (.A1(load),
    .A2(in_data_flat[67]),
    .B1(_0192_),
    .B2(\gen_left[2][3] ),
    .X(_2214_));
 sky130_fd_sc_hd__a21o_2 _2667_ (.A1(\gen_pe[1].pe_inst.out_right[3] ),
    .A2(_1543_),
    .B1(_2214_),
    .X(_0057_));
 sky130_fd_sc_hd__a22o_2 _2668_ (.A1(load),
    .A2(in_data_flat[68]),
    .B1(_0192_),
    .B2(\gen_left[2][4] ),
    .X(_2215_));
 sky130_fd_sc_hd__a21o_2 _2669_ (.A1(\gen_pe[1].pe_inst.out_right[4] ),
    .A2(_1543_),
    .B1(_2215_),
    .X(_0058_));
 sky130_fd_sc_hd__a22o_2 _2670_ (.A1(load),
    .A2(in_data_flat[69]),
    .B1(_0192_),
    .B2(\gen_left[2][5] ),
    .X(_2216_));
 sky130_fd_sc_hd__a21o_2 _2671_ (.A1(\gen_pe[1].pe_inst.out_right[5] ),
    .A2(_1543_),
    .B1(_2216_),
    .X(_0059_));
 sky130_fd_sc_hd__a22o_2 _2672_ (.A1(load),
    .A2(in_data_flat[70]),
    .B1(_0192_),
    .B2(\gen_left[2][6] ),
    .X(_2217_));
 sky130_fd_sc_hd__a21o_2 _2673_ (.A1(\gen_pe[1].pe_inst.out_right[6] ),
    .A2(_1543_),
    .B1(_2217_),
    .X(_0060_));
 sky130_fd_sc_hd__and2_2 _2674_ (.A(load),
    .B(in_data_flat[71]),
    .X(_2218_));
 sky130_fd_sc_hd__a221o_2 _2675_ (.A1(\gen_left[2][7] ),
    .A2(_0192_),
    .B1(_1543_),
    .B2(\gen_pe[1].pe_inst.out_right[7] ),
    .C1(_2218_),
    .X(_0061_));
 sky130_fd_sc_hd__a22o_2 _2676_ (.A1(load),
    .A2(in_data_flat[72]),
    .B1(_0192_),
    .B2(\gen_left[2][8] ),
    .X(_2219_));
 sky130_fd_sc_hd__a21o_2 _2677_ (.A1(\gen_pe[1].pe_inst.out_right[8] ),
    .A2(_1543_),
    .B1(_2219_),
    .X(_0062_));
 sky130_fd_sc_hd__a22o_2 _2678_ (.A1(load),
    .A2(in_data_flat[73]),
    .B1(_0192_),
    .B2(\gen_left[2][9] ),
    .X(_2220_));
 sky130_fd_sc_hd__a21o_2 _2679_ (.A1(\gen_pe[1].pe_inst.out_right[9] ),
    .A2(_1543_),
    .B1(_2220_),
    .X(_0063_));
 sky130_fd_sc_hd__a22o_2 _2680_ (.A1(load),
    .A2(in_data_flat[74]),
    .B1(_0192_),
    .B2(\gen_left[2][10] ),
    .X(_2221_));
 sky130_fd_sc_hd__a21o_2 _2681_ (.A1(\gen_pe[1].pe_inst.out_right[10] ),
    .A2(_1543_),
    .B1(_2221_),
    .X(_0033_));
 sky130_fd_sc_hd__a22o_2 _2682_ (.A1(load),
    .A2(in_data_flat[75]),
    .B1(_0192_),
    .B2(\gen_left[2][11] ),
    .X(_2222_));
 sky130_fd_sc_hd__a21o_2 _2683_ (.A1(\gen_pe[1].pe_inst.out_right[11] ),
    .A2(_1543_),
    .B1(_2222_),
    .X(_0034_));
 sky130_fd_sc_hd__a22o_2 _2684_ (.A1(load),
    .A2(in_data_flat[76]),
    .B1(_0192_),
    .B2(\gen_left[2][12] ),
    .X(_2223_));
 sky130_fd_sc_hd__a21o_2 _2685_ (.A1(\gen_pe[1].pe_inst.out_right[12] ),
    .A2(_1543_),
    .B1(_2223_),
    .X(_0035_));
 sky130_fd_sc_hd__a22o_2 _2686_ (.A1(load),
    .A2(in_data_flat[77]),
    .B1(_0192_),
    .B2(\gen_left[2][13] ),
    .X(_2224_));
 sky130_fd_sc_hd__a21o_2 _2687_ (.A1(\gen_pe[1].pe_inst.out_right[13] ),
    .A2(_1543_),
    .B1(_2224_),
    .X(_0036_));
 sky130_fd_sc_hd__and2_2 _2688_ (.A(load),
    .B(in_data_flat[78]),
    .X(_2225_));
 sky130_fd_sc_hd__a221o_2 _2689_ (.A1(\gen_left[2][14] ),
    .A2(_0192_),
    .B1(_1543_),
    .B2(\gen_pe[1].pe_inst.out_right[14] ),
    .C1(_2225_),
    .X(_0037_));
 sky130_fd_sc_hd__and2_2 _2690_ (.A(load),
    .B(in_data_flat[79]),
    .X(_2226_));
 sky130_fd_sc_hd__a221o_2 _2691_ (.A1(\gen_left[2][15] ),
    .A2(_0192_),
    .B1(_1543_),
    .B2(\gen_pe[1].pe_inst.out_right[15] ),
    .C1(_2226_),
    .X(_0038_));
 sky130_fd_sc_hd__a22o_2 _2692_ (.A1(load),
    .A2(in_data_flat[80]),
    .B1(_0192_),
    .B2(\gen_left[2][16] ),
    .X(_2227_));
 sky130_fd_sc_hd__a21o_2 _2693_ (.A1(\gen_pe[1].pe_inst.out_right[16] ),
    .A2(_1543_),
    .B1(_2227_),
    .X(_0039_));
 sky130_fd_sc_hd__a22o_2 _2694_ (.A1(load),
    .A2(in_data_flat[81]),
    .B1(_0192_),
    .B2(\gen_left[2][17] ),
    .X(_2228_));
 sky130_fd_sc_hd__a21o_2 _2695_ (.A1(\gen_pe[1].pe_inst.out_right[17] ),
    .A2(_1543_),
    .B1(_2228_),
    .X(_0040_));
 sky130_fd_sc_hd__a22o_2 _2696_ (.A1(load),
    .A2(in_data_flat[82]),
    .B1(_0192_),
    .B2(\gen_left[2][18] ),
    .X(_2229_));
 sky130_fd_sc_hd__a21o_2 _2697_ (.A1(\gen_pe[1].pe_inst.out_right[18] ),
    .A2(_1543_),
    .B1(_2229_),
    .X(_0041_));
 sky130_fd_sc_hd__a22o_2 _2698_ (.A1(load),
    .A2(in_data_flat[83]),
    .B1(_0192_),
    .B2(\gen_left[2][19] ),
    .X(_2230_));
 sky130_fd_sc_hd__a21o_2 _2699_ (.A1(\gen_pe[1].pe_inst.out_right[19] ),
    .A2(_1543_),
    .B1(_2230_),
    .X(_0042_));
 sky130_fd_sc_hd__a22o_2 _2700_ (.A1(load),
    .A2(in_data_flat[84]),
    .B1(_0192_),
    .B2(\gen_left[2][20] ),
    .X(_2231_));
 sky130_fd_sc_hd__a21o_2 _2701_ (.A1(\gen_pe[1].pe_inst.out_right[20] ),
    .A2(_1543_),
    .B1(_2231_),
    .X(_0044_));
 sky130_fd_sc_hd__a22o_2 _2702_ (.A1(load),
    .A2(in_data_flat[85]),
    .B1(_0192_),
    .B2(\gen_left[2][21] ),
    .X(_2232_));
 sky130_fd_sc_hd__a21o_2 _2703_ (.A1(\gen_pe[1].pe_inst.out_right[21] ),
    .A2(_1543_),
    .B1(_2232_),
    .X(_0045_));
 sky130_fd_sc_hd__a22o_2 _2704_ (.A1(load),
    .A2(in_data_flat[86]),
    .B1(_0192_),
    .B2(\gen_left[2][22] ),
    .X(_2233_));
 sky130_fd_sc_hd__a21o_2 _2705_ (.A1(\gen_pe[1].pe_inst.out_right[22] ),
    .A2(_1543_),
    .B1(_2233_),
    .X(_0046_));
 sky130_fd_sc_hd__a22o_2 _2706_ (.A1(load),
    .A2(in_data_flat[87]),
    .B1(_0192_),
    .B2(\gen_left[2][23] ),
    .X(_2234_));
 sky130_fd_sc_hd__a21o_2 _2707_ (.A1(\gen_pe[1].pe_inst.out_right[23] ),
    .A2(_1543_),
    .B1(_2234_),
    .X(_0047_));
 sky130_fd_sc_hd__a22o_2 _2708_ (.A1(load),
    .A2(in_data_flat[88]),
    .B1(_0192_),
    .B2(\gen_left[2][24] ),
    .X(_2235_));
 sky130_fd_sc_hd__a21o_2 _2709_ (.A1(\gen_pe[1].pe_inst.out_right[24] ),
    .A2(_1543_),
    .B1(_2235_),
    .X(_0048_));
 sky130_fd_sc_hd__and2_2 _2710_ (.A(load),
    .B(in_data_flat[89]),
    .X(_2236_));
 sky130_fd_sc_hd__a221o_2 _2711_ (.A1(\gen_left[2][25] ),
    .A2(_0192_),
    .B1(_1543_),
    .B2(\gen_pe[1].pe_inst.out_right[25] ),
    .C1(_2236_),
    .X(_0049_));
 sky130_fd_sc_hd__a22o_2 _2712_ (.A1(load),
    .A2(in_data_flat[90]),
    .B1(_0192_),
    .B2(\gen_left[2][26] ),
    .X(_2237_));
 sky130_fd_sc_hd__a21o_2 _2713_ (.A1(\gen_pe[1].pe_inst.out_right[26] ),
    .A2(_1543_),
    .B1(_2237_),
    .X(_0050_));
 sky130_fd_sc_hd__a22o_2 _2714_ (.A1(load),
    .A2(in_data_flat[91]),
    .B1(_0192_),
    .B2(\gen_left[2][27] ),
    .X(_2238_));
 sky130_fd_sc_hd__a21o_2 _2715_ (.A1(\gen_pe[1].pe_inst.out_right[27] ),
    .A2(_1543_),
    .B1(_2238_),
    .X(_0051_));
 sky130_fd_sc_hd__and2_2 _2716_ (.A(load),
    .B(in_data_flat[92]),
    .X(_2239_));
 sky130_fd_sc_hd__a221o_2 _2717_ (.A1(\gen_left[2][28] ),
    .A2(_0192_),
    .B1(_1543_),
    .B2(\gen_pe[1].pe_inst.out_right[28] ),
    .C1(_2239_),
    .X(_0052_));
 sky130_fd_sc_hd__a22o_2 _2718_ (.A1(load),
    .A2(in_data_flat[93]),
    .B1(_0192_),
    .B2(\gen_left[2][29] ),
    .X(_2240_));
 sky130_fd_sc_hd__a21o_2 _2719_ (.A1(\gen_pe[1].pe_inst.out_right[29] ),
    .A2(_1543_),
    .B1(_2240_),
    .X(_0053_));
 sky130_fd_sc_hd__a22o_2 _2720_ (.A1(load),
    .A2(in_data_flat[94]),
    .B1(_0192_),
    .B2(\gen_left[2][30] ),
    .X(_2241_));
 sky130_fd_sc_hd__a21o_2 _2721_ (.A1(\gen_pe[1].pe_inst.out_right[30] ),
    .A2(_1543_),
    .B1(_2241_),
    .X(_0055_));
 sky130_fd_sc_hd__a22o_2 _2722_ (.A1(load),
    .A2(in_data_flat[95]),
    .B1(_0192_),
    .B2(\gen_left[2][31] ),
    .X(_2242_));
 sky130_fd_sc_hd__a21o_2 _2723_ (.A1(\gen_pe[1].pe_inst.out_right[31] ),
    .A2(_1543_),
    .B1(_2242_),
    .X(_0056_));
 sky130_fd_sc_hd__a22o_2 _2724_ (.A1(load),
    .A2(in_data_flat[96]),
    .B1(_0192_),
    .B2(\gen_pe[2].pe_inst.out_right[0] ),
    .X(_2243_));
 sky130_fd_sc_hd__a21o_2 _2725_ (.A1(\gen_left[3][0] ),
    .A2(_1543_),
    .B1(_2243_),
    .X(_0064_));
 sky130_fd_sc_hd__a22o_2 _2726_ (.A1(load),
    .A2(in_data_flat[97]),
    .B1(_0192_),
    .B2(\gen_pe[2].pe_inst.out_right[1] ),
    .X(_2244_));
 sky130_fd_sc_hd__a21o_2 _2727_ (.A1(\gen_left[3][1] ),
    .A2(_1543_),
    .B1(_2244_),
    .X(_0075_));
 sky130_fd_sc_hd__a22o_2 _2728_ (.A1(load),
    .A2(in_data_flat[98]),
    .B1(_0192_),
    .B2(\gen_pe[2].pe_inst.out_right[2] ),
    .X(_2245_));
 sky130_fd_sc_hd__a21o_2 _2729_ (.A1(\gen_left[3][2] ),
    .A2(_1543_),
    .B1(_2245_),
    .X(_0086_));
 sky130_fd_sc_hd__a22o_2 _2730_ (.A1(load),
    .A2(in_data_flat[99]),
    .B1(_0192_),
    .B2(\gen_pe[2].pe_inst.out_right[3] ),
    .X(_2246_));
 sky130_fd_sc_hd__a21o_2 _2731_ (.A1(\gen_left[3][3] ),
    .A2(_1543_),
    .B1(_2246_),
    .X(_0089_));
 sky130_fd_sc_hd__a22o_2 _2732_ (.A1(load),
    .A2(in_data_flat[100]),
    .B1(_0192_),
    .B2(\gen_pe[2].pe_inst.out_right[4] ),
    .X(_2247_));
 sky130_fd_sc_hd__a21o_2 _2733_ (.A1(\gen_left[3][4] ),
    .A2(_1543_),
    .B1(_2247_),
    .X(_0090_));
 sky130_fd_sc_hd__a22o_2 _2734_ (.A1(load),
    .A2(in_data_flat[101]),
    .B1(_0192_),
    .B2(\gen_pe[2].pe_inst.out_right[5] ),
    .X(_2248_));
 sky130_fd_sc_hd__a21o_2 _2735_ (.A1(\gen_left[3][5] ),
    .A2(_1543_),
    .B1(_2248_),
    .X(_0091_));
 sky130_fd_sc_hd__a22o_2 _2736_ (.A1(load),
    .A2(in_data_flat[102]),
    .B1(_0192_),
    .B2(\gen_pe[2].pe_inst.out_right[6] ),
    .X(_2249_));
 sky130_fd_sc_hd__a21o_2 _2737_ (.A1(\gen_left[3][6] ),
    .A2(_1543_),
    .B1(_2249_),
    .X(_0092_));
 sky130_fd_sc_hd__and2_2 _2738_ (.A(load),
    .B(in_data_flat[103]),
    .X(_2250_));
 sky130_fd_sc_hd__a221o_2 _2739_ (.A1(\gen_pe[2].pe_inst.out_right[7] ),
    .A2(_0192_),
    .B1(_1543_),
    .B2(\gen_left[3][7] ),
    .C1(_2250_),
    .X(_0093_));
 sky130_fd_sc_hd__a22o_2 _2740_ (.A1(load),
    .A2(in_data_flat[104]),
    .B1(_0192_),
    .B2(\gen_pe[2].pe_inst.out_right[8] ),
    .X(_2251_));
 sky130_fd_sc_hd__a21o_2 _2741_ (.A1(\gen_left[3][8] ),
    .A2(_1543_),
    .B1(_2251_),
    .X(_0094_));
 sky130_fd_sc_hd__a22o_2 _2742_ (.A1(load),
    .A2(in_data_flat[105]),
    .B1(_0192_),
    .B2(\gen_pe[2].pe_inst.out_right[9] ),
    .X(_2252_));
 sky130_fd_sc_hd__a21o_2 _2743_ (.A1(\gen_left[3][9] ),
    .A2(_1543_),
    .B1(_2252_),
    .X(_0095_));
 sky130_fd_sc_hd__a22o_2 _2744_ (.A1(load),
    .A2(in_data_flat[106]),
    .B1(_0192_),
    .B2(\gen_pe[2].pe_inst.out_right[10] ),
    .X(_2253_));
 sky130_fd_sc_hd__a21o_2 _2745_ (.A1(\gen_left[3][10] ),
    .A2(_1543_),
    .B1(_2253_),
    .X(_0065_));
 sky130_fd_sc_hd__a22o_2 _2746_ (.A1(load),
    .A2(in_data_flat[107]),
    .B1(_0192_),
    .B2(\gen_pe[2].pe_inst.out_right[11] ),
    .X(_2254_));
 sky130_fd_sc_hd__a21o_2 _2747_ (.A1(\gen_left[3][11] ),
    .A2(_1543_),
    .B1(_2254_),
    .X(_0066_));
 sky130_fd_sc_hd__a22o_2 _2748_ (.A1(load),
    .A2(in_data_flat[108]),
    .B1(_0192_),
    .B2(\gen_pe[2].pe_inst.out_right[12] ),
    .X(_2255_));
 sky130_fd_sc_hd__a21o_2 _2749_ (.A1(\gen_left[3][12] ),
    .A2(_1543_),
    .B1(_2255_),
    .X(_0067_));
 sky130_fd_sc_hd__a22o_2 _2750_ (.A1(load),
    .A2(in_data_flat[109]),
    .B1(_0192_),
    .B2(\gen_pe[2].pe_inst.out_right[13] ),
    .X(_2256_));
 sky130_fd_sc_hd__a21o_2 _2751_ (.A1(\gen_left[3][13] ),
    .A2(_1543_),
    .B1(_2256_),
    .X(_0068_));
 sky130_fd_sc_hd__and2_2 _2752_ (.A(load),
    .B(in_data_flat[110]),
    .X(_2257_));
 sky130_fd_sc_hd__a221o_2 _2753_ (.A1(\gen_pe[2].pe_inst.out_right[14] ),
    .A2(_0192_),
    .B1(_1543_),
    .B2(\gen_left[3][14] ),
    .C1(_2257_),
    .X(_0069_));
 sky130_fd_sc_hd__and2_2 _2754_ (.A(load),
    .B(in_data_flat[111]),
    .X(_2258_));
 sky130_fd_sc_hd__a221o_2 _2755_ (.A1(\gen_pe[2].pe_inst.out_right[15] ),
    .A2(_0192_),
    .B1(_1543_),
    .B2(\gen_left[3][15] ),
    .C1(_2258_),
    .X(_0070_));
 sky130_fd_sc_hd__a22o_2 _2756_ (.A1(load),
    .A2(in_data_flat[112]),
    .B1(_0192_),
    .B2(\gen_pe[2].pe_inst.out_right[16] ),
    .X(_2259_));
 sky130_fd_sc_hd__a21o_2 _2757_ (.A1(\gen_left[3][16] ),
    .A2(_1543_),
    .B1(_2259_),
    .X(_0071_));
 sky130_fd_sc_hd__a22o_2 _2758_ (.A1(load),
    .A2(in_data_flat[113]),
    .B1(_0192_),
    .B2(\gen_pe[2].pe_inst.out_right[17] ),
    .X(_2260_));
 sky130_fd_sc_hd__a21o_2 _2759_ (.A1(\gen_left[3][17] ),
    .A2(_1543_),
    .B1(_2260_),
    .X(_0072_));
 sky130_fd_sc_hd__a22o_2 _2760_ (.A1(load),
    .A2(in_data_flat[114]),
    .B1(_0192_),
    .B2(\gen_pe[2].pe_inst.out_right[18] ),
    .X(_2261_));
 sky130_fd_sc_hd__a21o_2 _2761_ (.A1(\gen_left[3][18] ),
    .A2(_1543_),
    .B1(_2261_),
    .X(_0073_));
 sky130_fd_sc_hd__a22o_2 _2762_ (.A1(load),
    .A2(in_data_flat[115]),
    .B1(_0192_),
    .B2(\gen_pe[2].pe_inst.out_right[19] ),
    .X(_2262_));
 sky130_fd_sc_hd__a21o_2 _2763_ (.A1(\gen_left[3][19] ),
    .A2(_1543_),
    .B1(_2262_),
    .X(_0074_));
 sky130_fd_sc_hd__a22o_2 _2764_ (.A1(load),
    .A2(in_data_flat[116]),
    .B1(_0192_),
    .B2(\gen_pe[2].pe_inst.out_right[20] ),
    .X(_2263_));
 sky130_fd_sc_hd__a21o_2 _2765_ (.A1(\gen_left[3][20] ),
    .A2(_1543_),
    .B1(_2263_),
    .X(_0076_));
 sky130_fd_sc_hd__a22o_2 _2766_ (.A1(load),
    .A2(in_data_flat[117]),
    .B1(_0192_),
    .B2(\gen_pe[2].pe_inst.out_right[21] ),
    .X(_2264_));
 sky130_fd_sc_hd__a21o_2 _2767_ (.A1(\gen_left[3][21] ),
    .A2(_1543_),
    .B1(_2264_),
    .X(_0077_));
 sky130_fd_sc_hd__a22o_2 _2768_ (.A1(load),
    .A2(in_data_flat[118]),
    .B1(_0192_),
    .B2(\gen_pe[2].pe_inst.out_right[22] ),
    .X(_2265_));
 sky130_fd_sc_hd__a21o_2 _2769_ (.A1(\gen_left[3][22] ),
    .A2(_1543_),
    .B1(_2265_),
    .X(_0078_));
 sky130_fd_sc_hd__a22o_2 _2770_ (.A1(load),
    .A2(in_data_flat[119]),
    .B1(_0192_),
    .B2(\gen_pe[2].pe_inst.out_right[23] ),
    .X(_2266_));
 sky130_fd_sc_hd__a21o_2 _2771_ (.A1(\gen_left[3][23] ),
    .A2(_1543_),
    .B1(_2266_),
    .X(_0079_));
 sky130_fd_sc_hd__a22o_2 _2772_ (.A1(load),
    .A2(in_data_flat[120]),
    .B1(_0192_),
    .B2(\gen_pe[2].pe_inst.out_right[24] ),
    .X(_2267_));
 sky130_fd_sc_hd__a21o_2 _2773_ (.A1(\gen_left[3][24] ),
    .A2(_1543_),
    .B1(_2267_),
    .X(_0080_));
 sky130_fd_sc_hd__and2_2 _2774_ (.A(load),
    .B(in_data_flat[121]),
    .X(_2268_));
 sky130_fd_sc_hd__a221o_2 _2775_ (.A1(\gen_pe[2].pe_inst.out_right[25] ),
    .A2(_0192_),
    .B1(_1543_),
    .B2(\gen_left[3][25] ),
    .C1(_2268_),
    .X(_0081_));
 sky130_fd_sc_hd__a22o_2 _2776_ (.A1(load),
    .A2(in_data_flat[122]),
    .B1(_0192_),
    .B2(\gen_pe[2].pe_inst.out_right[26] ),
    .X(_2269_));
 sky130_fd_sc_hd__a21o_2 _2777_ (.A1(\gen_left[3][26] ),
    .A2(_1543_),
    .B1(_2269_),
    .X(_0082_));
 sky130_fd_sc_hd__a22o_2 _2778_ (.A1(load),
    .A2(in_data_flat[123]),
    .B1(_0192_),
    .B2(\gen_pe[2].pe_inst.out_right[27] ),
    .X(_2270_));
 sky130_fd_sc_hd__a21o_2 _2779_ (.A1(\gen_left[3][27] ),
    .A2(_1543_),
    .B1(_2270_),
    .X(_0083_));
 sky130_fd_sc_hd__and2_2 _2780_ (.A(load),
    .B(in_data_flat[124]),
    .X(_2271_));
 sky130_fd_sc_hd__a221o_2 _2781_ (.A1(\gen_pe[2].pe_inst.out_right[28] ),
    .A2(_0192_),
    .B1(_1543_),
    .B2(\gen_left[3][28] ),
    .C1(_2271_),
    .X(_0084_));
 sky130_fd_sc_hd__a22o_2 _2782_ (.A1(load),
    .A2(in_data_flat[125]),
    .B1(_0192_),
    .B2(\gen_pe[2].pe_inst.out_right[29] ),
    .X(_2272_));
 sky130_fd_sc_hd__a21o_2 _2783_ (.A1(\gen_left[3][29] ),
    .A2(_1543_),
    .B1(_2272_),
    .X(_0085_));
 sky130_fd_sc_hd__a22o_2 _2784_ (.A1(load),
    .A2(in_data_flat[126]),
    .B1(_0192_),
    .B2(\gen_pe[2].pe_inst.out_right[30] ),
    .X(_2273_));
 sky130_fd_sc_hd__a21o_2 _2785_ (.A1(\gen_left[3][30] ),
    .A2(_1543_),
    .B1(_2273_),
    .X(_0087_));
 sky130_fd_sc_hd__a22o_2 _2786_ (.A1(load),
    .A2(in_data_flat[127]),
    .B1(_0192_),
    .B2(\gen_pe[2].pe_inst.out_right[31] ),
    .X(_2274_));
 sky130_fd_sc_hd__a21o_2 _2787_ (.A1(\gen_left[3][31] ),
    .A2(_1543_),
    .B1(_2274_),
    .X(_0088_));
 sky130_fd_sc_hd__a22o_2 _2788_ (.A1(load),
    .A2(in_data_flat[128]),
    .B1(_0192_),
    .B2(\gen_left[4][0] ),
    .X(_2275_));
 sky130_fd_sc_hd__a21o_2 _2789_ (.A1(\gen_pe[3].pe_inst.out_right[0] ),
    .A2(_1543_),
    .B1(_2275_),
    .X(_0096_));
 sky130_fd_sc_hd__a22o_2 _2790_ (.A1(load),
    .A2(in_data_flat[129]),
    .B1(_0192_),
    .B2(\gen_left[4][1] ),
    .X(_2276_));
 sky130_fd_sc_hd__a21o_2 _2791_ (.A1(\gen_pe[3].pe_inst.out_right[1] ),
    .A2(_1543_),
    .B1(_2276_),
    .X(_0107_));
 sky130_fd_sc_hd__a22o_2 _2792_ (.A1(load),
    .A2(in_data_flat[130]),
    .B1(_0192_),
    .B2(\gen_left[4][2] ),
    .X(_2277_));
 sky130_fd_sc_hd__a21o_2 _2793_ (.A1(\gen_pe[3].pe_inst.out_right[2] ),
    .A2(_1543_),
    .B1(_2277_),
    .X(_0118_));
 sky130_fd_sc_hd__a22o_2 _2794_ (.A1(load),
    .A2(in_data_flat[131]),
    .B1(_0192_),
    .B2(\gen_left[4][3] ),
    .X(_2278_));
 sky130_fd_sc_hd__a21o_2 _2795_ (.A1(\gen_pe[3].pe_inst.out_right[3] ),
    .A2(_1543_),
    .B1(_2278_),
    .X(_0121_));
 sky130_fd_sc_hd__a22o_2 _2796_ (.A1(load),
    .A2(in_data_flat[132]),
    .B1(_0192_),
    .B2(\gen_left[4][4] ),
    .X(_2279_));
 sky130_fd_sc_hd__a21o_2 _2797_ (.A1(\gen_pe[3].pe_inst.out_right[4] ),
    .A2(_1543_),
    .B1(_2279_),
    .X(_0122_));
 sky130_fd_sc_hd__a22o_2 _2798_ (.A1(load),
    .A2(in_data_flat[133]),
    .B1(_0192_),
    .B2(\gen_left[4][5] ),
    .X(_2280_));
 sky130_fd_sc_hd__a21o_2 _2799_ (.A1(\gen_pe[3].pe_inst.out_right[5] ),
    .A2(_1543_),
    .B1(_2280_),
    .X(_0123_));
 sky130_fd_sc_hd__a22o_2 _2800_ (.A1(load),
    .A2(in_data_flat[134]),
    .B1(_0192_),
    .B2(\gen_left[4][6] ),
    .X(_2281_));
 sky130_fd_sc_hd__a21o_2 _2801_ (.A1(\gen_pe[3].pe_inst.out_right[6] ),
    .A2(_1543_),
    .B1(_2281_),
    .X(_0124_));
 sky130_fd_sc_hd__and2_2 _2802_ (.A(load),
    .B(in_data_flat[135]),
    .X(_2282_));
 sky130_fd_sc_hd__a221o_2 _2803_ (.A1(\gen_left[4][7] ),
    .A2(_0192_),
    .B1(_1543_),
    .B2(\gen_pe[3].pe_inst.out_right[7] ),
    .C1(_2282_),
    .X(_0125_));
 sky130_fd_sc_hd__a22o_2 _2804_ (.A1(load),
    .A2(in_data_flat[136]),
    .B1(_0192_),
    .B2(\gen_left[4][8] ),
    .X(_2283_));
 sky130_fd_sc_hd__a21o_2 _2805_ (.A1(\gen_pe[3].pe_inst.out_right[8] ),
    .A2(_1543_),
    .B1(_2283_),
    .X(_0126_));
 sky130_fd_sc_hd__a22o_2 _2806_ (.A1(load),
    .A2(in_data_flat[137]),
    .B1(_0192_),
    .B2(\gen_left[4][9] ),
    .X(_2284_));
 sky130_fd_sc_hd__a21o_2 _2807_ (.A1(\gen_pe[3].pe_inst.out_right[9] ),
    .A2(_1543_),
    .B1(_2284_),
    .X(_0127_));
 sky130_fd_sc_hd__a22o_2 _2808_ (.A1(load),
    .A2(in_data_flat[138]),
    .B1(_0192_),
    .B2(\gen_left[4][10] ),
    .X(_2285_));
 sky130_fd_sc_hd__a21o_2 _2809_ (.A1(\gen_pe[3].pe_inst.out_right[10] ),
    .A2(_1543_),
    .B1(_2285_),
    .X(_0097_));
 sky130_fd_sc_hd__a22o_2 _2810_ (.A1(load),
    .A2(in_data_flat[139]),
    .B1(_0192_),
    .B2(\gen_left[4][11] ),
    .X(_2286_));
 sky130_fd_sc_hd__a21o_2 _2811_ (.A1(\gen_pe[3].pe_inst.out_right[11] ),
    .A2(_1543_),
    .B1(_2286_),
    .X(_0098_));
 sky130_fd_sc_hd__a22o_2 _2812_ (.A1(load),
    .A2(in_data_flat[140]),
    .B1(_0192_),
    .B2(\gen_left[4][12] ),
    .X(_2287_));
 sky130_fd_sc_hd__a21o_2 _2813_ (.A1(\gen_pe[3].pe_inst.out_right[12] ),
    .A2(_1543_),
    .B1(_2287_),
    .X(_0099_));
 sky130_fd_sc_hd__a22o_2 _2814_ (.A1(load),
    .A2(in_data_flat[141]),
    .B1(_0192_),
    .B2(\gen_left[4][13] ),
    .X(_2288_));
 sky130_fd_sc_hd__a21o_2 _2815_ (.A1(\gen_pe[3].pe_inst.out_right[13] ),
    .A2(_1543_),
    .B1(_2288_),
    .X(_0100_));
 sky130_fd_sc_hd__and2_2 _2816_ (.A(load),
    .B(in_data_flat[142]),
    .X(_2289_));
 sky130_fd_sc_hd__a221o_2 _2817_ (.A1(\gen_left[4][14] ),
    .A2(_0192_),
    .B1(_1543_),
    .B2(\gen_pe[3].pe_inst.out_right[14] ),
    .C1(_2289_),
    .X(_0101_));
 sky130_fd_sc_hd__and2_2 _2818_ (.A(load),
    .B(in_data_flat[143]),
    .X(_2290_));
 sky130_fd_sc_hd__a221o_2 _2819_ (.A1(\gen_left[4][15] ),
    .A2(_0192_),
    .B1(_1543_),
    .B2(\gen_pe[3].pe_inst.out_right[15] ),
    .C1(_2290_),
    .X(_0102_));
 sky130_fd_sc_hd__a22o_2 _2820_ (.A1(load),
    .A2(in_data_flat[144]),
    .B1(_0192_),
    .B2(\gen_left[4][16] ),
    .X(_2291_));
 sky130_fd_sc_hd__a21o_2 _2821_ (.A1(\gen_pe[3].pe_inst.out_right[16] ),
    .A2(_1543_),
    .B1(_2291_),
    .X(_0103_));
 sky130_fd_sc_hd__a22o_2 _2822_ (.A1(load),
    .A2(in_data_flat[145]),
    .B1(_0192_),
    .B2(\gen_left[4][17] ),
    .X(_2292_));
 sky130_fd_sc_hd__a21o_2 _2823_ (.A1(\gen_pe[3].pe_inst.out_right[17] ),
    .A2(_1543_),
    .B1(_2292_),
    .X(_0104_));
 sky130_fd_sc_hd__a22o_2 _2824_ (.A1(load),
    .A2(in_data_flat[146]),
    .B1(_0192_),
    .B2(\gen_left[4][18] ),
    .X(_2293_));
 sky130_fd_sc_hd__a21o_2 _2825_ (.A1(\gen_pe[3].pe_inst.out_right[18] ),
    .A2(_1543_),
    .B1(_2293_),
    .X(_0105_));
 sky130_fd_sc_hd__a22o_2 _2826_ (.A1(load),
    .A2(in_data_flat[147]),
    .B1(_0192_),
    .B2(\gen_left[4][19] ),
    .X(_2294_));
 sky130_fd_sc_hd__a21o_2 _2827_ (.A1(\gen_pe[3].pe_inst.out_right[19] ),
    .A2(_1543_),
    .B1(_2294_),
    .X(_0106_));
 sky130_fd_sc_hd__a22o_2 _2828_ (.A1(load),
    .A2(in_data_flat[148]),
    .B1(_0192_),
    .B2(\gen_left[4][20] ),
    .X(_2295_));
 sky130_fd_sc_hd__a21o_2 _2829_ (.A1(\gen_pe[3].pe_inst.out_right[20] ),
    .A2(_1543_),
    .B1(_2295_),
    .X(_0108_));
 sky130_fd_sc_hd__a22o_2 _2830_ (.A1(load),
    .A2(in_data_flat[149]),
    .B1(_0192_),
    .B2(\gen_left[4][21] ),
    .X(_2296_));
 sky130_fd_sc_hd__a21o_2 _2831_ (.A1(\gen_pe[3].pe_inst.out_right[21] ),
    .A2(_1543_),
    .B1(_2296_),
    .X(_0109_));
 sky130_fd_sc_hd__a22o_2 _2832_ (.A1(load),
    .A2(in_data_flat[150]),
    .B1(_0192_),
    .B2(\gen_left[4][22] ),
    .X(_2297_));
 sky130_fd_sc_hd__a21o_2 _2833_ (.A1(\gen_pe[3].pe_inst.out_right[22] ),
    .A2(_1543_),
    .B1(_2297_),
    .X(_0110_));
 sky130_fd_sc_hd__a22o_2 _2834_ (.A1(load),
    .A2(in_data_flat[151]),
    .B1(_0192_),
    .B2(\gen_left[4][23] ),
    .X(_2298_));
 sky130_fd_sc_hd__a21o_2 _2835_ (.A1(\gen_pe[3].pe_inst.out_right[23] ),
    .A2(_1543_),
    .B1(_2298_),
    .X(_0111_));
 sky130_fd_sc_hd__a22o_2 _2836_ (.A1(load),
    .A2(in_data_flat[152]),
    .B1(_0192_),
    .B2(\gen_left[4][24] ),
    .X(_2299_));
 sky130_fd_sc_hd__a21o_2 _2837_ (.A1(\gen_pe[3].pe_inst.out_right[24] ),
    .A2(_1543_),
    .B1(_2299_),
    .X(_0112_));
 sky130_fd_sc_hd__and2_2 _2838_ (.A(load),
    .B(in_data_flat[153]),
    .X(_2300_));
 sky130_fd_sc_hd__a221o_2 _2839_ (.A1(\gen_left[4][25] ),
    .A2(_0192_),
    .B1(_1543_),
    .B2(\gen_pe[3].pe_inst.out_right[25] ),
    .C1(_2300_),
    .X(_0113_));
 sky130_fd_sc_hd__a22o_2 _2840_ (.A1(load),
    .A2(in_data_flat[154]),
    .B1(_0192_),
    .B2(\gen_left[4][26] ),
    .X(_2301_));
 sky130_fd_sc_hd__a21o_2 _2841_ (.A1(\gen_pe[3].pe_inst.out_right[26] ),
    .A2(_1543_),
    .B1(_2301_),
    .X(_0114_));
 sky130_fd_sc_hd__a22o_2 _2842_ (.A1(load),
    .A2(in_data_flat[155]),
    .B1(_0192_),
    .B2(\gen_left[4][27] ),
    .X(_2302_));
 sky130_fd_sc_hd__a21o_2 _2843_ (.A1(\gen_pe[3].pe_inst.out_right[27] ),
    .A2(_1543_),
    .B1(_2302_),
    .X(_0115_));
 sky130_fd_sc_hd__and2_2 _2844_ (.A(load),
    .B(in_data_flat[156]),
    .X(_2303_));
 sky130_fd_sc_hd__a221o_2 _2845_ (.A1(\gen_left[4][28] ),
    .A2(_0192_),
    .B1(_1543_),
    .B2(\gen_pe[3].pe_inst.out_right[28] ),
    .C1(_2303_),
    .X(_0116_));
 sky130_fd_sc_hd__a22o_2 _2846_ (.A1(load),
    .A2(in_data_flat[157]),
    .B1(_0192_),
    .B2(\gen_left[4][29] ),
    .X(_2304_));
 sky130_fd_sc_hd__a21o_2 _2847_ (.A1(\gen_pe[3].pe_inst.out_right[29] ),
    .A2(_1543_),
    .B1(_2304_),
    .X(_0117_));
 sky130_fd_sc_hd__a22o_2 _2848_ (.A1(load),
    .A2(in_data_flat[158]),
    .B1(_0192_),
    .B2(\gen_left[4][30] ),
    .X(_2305_));
 sky130_fd_sc_hd__a21o_2 _2849_ (.A1(\gen_pe[3].pe_inst.out_right[30] ),
    .A2(_1543_),
    .B1(_2305_),
    .X(_0119_));
 sky130_fd_sc_hd__a22o_2 _2850_ (.A1(load),
    .A2(in_data_flat[159]),
    .B1(_0192_),
    .B2(\gen_left[4][31] ),
    .X(_2306_));
 sky130_fd_sc_hd__a21o_2 _2851_ (.A1(\gen_pe[3].pe_inst.out_right[31] ),
    .A2(_1543_),
    .B1(_2306_),
    .X(_0120_));
 sky130_fd_sc_hd__a22o_2 _2852_ (.A1(load),
    .A2(in_data_flat[160]),
    .B1(_0192_),
    .B2(\gen_pe[4].pe_inst.out_right[0] ),
    .X(_2307_));
 sky130_fd_sc_hd__a21o_2 _2853_ (.A1(\gen_left[5][0] ),
    .A2(_1543_),
    .B1(_2307_),
    .X(_0128_));
 sky130_fd_sc_hd__a22o_2 _2854_ (.A1(load),
    .A2(in_data_flat[161]),
    .B1(_0192_),
    .B2(\gen_pe[4].pe_inst.out_right[1] ),
    .X(_2308_));
 sky130_fd_sc_hd__a21o_2 _2855_ (.A1(\gen_left[5][1] ),
    .A2(_1543_),
    .B1(_2308_),
    .X(_0139_));
 sky130_fd_sc_hd__a22o_2 _2856_ (.A1(load),
    .A2(in_data_flat[162]),
    .B1(_0192_),
    .B2(\gen_pe[4].pe_inst.out_right[2] ),
    .X(_2309_));
 sky130_fd_sc_hd__a21o_2 _2857_ (.A1(\gen_left[5][2] ),
    .A2(_1543_),
    .B1(_2309_),
    .X(_0150_));
 sky130_fd_sc_hd__a22o_2 _2858_ (.A1(load),
    .A2(in_data_flat[163]),
    .B1(_0192_),
    .B2(\gen_pe[4].pe_inst.out_right[3] ),
    .X(_2310_));
 sky130_fd_sc_hd__a21o_2 _2859_ (.A1(\gen_left[5][3] ),
    .A2(_1543_),
    .B1(_2310_),
    .X(_0153_));
 sky130_fd_sc_hd__a22o_2 _2860_ (.A1(load),
    .A2(in_data_flat[164]),
    .B1(_0192_),
    .B2(\gen_pe[4].pe_inst.out_right[4] ),
    .X(_2311_));
 sky130_fd_sc_hd__a21o_2 _2861_ (.A1(\gen_left[5][4] ),
    .A2(_1543_),
    .B1(_2311_),
    .X(_0154_));
 sky130_fd_sc_hd__a22o_2 _2862_ (.A1(load),
    .A2(in_data_flat[165]),
    .B1(_0192_),
    .B2(\gen_pe[4].pe_inst.out_right[5] ),
    .X(_2312_));
 sky130_fd_sc_hd__a21o_2 _2863_ (.A1(\gen_left[5][5] ),
    .A2(_1543_),
    .B1(_2312_),
    .X(_0155_));
 sky130_fd_sc_hd__a22o_2 _2864_ (.A1(load),
    .A2(in_data_flat[166]),
    .B1(_0192_),
    .B2(\gen_pe[4].pe_inst.out_right[6] ),
    .X(_2313_));
 sky130_fd_sc_hd__a21o_2 _2865_ (.A1(\gen_left[5][6] ),
    .A2(_1543_),
    .B1(_2313_),
    .X(_0156_));
 sky130_fd_sc_hd__and2_2 _2866_ (.A(load),
    .B(in_data_flat[167]),
    .X(_2314_));
 sky130_fd_sc_hd__a221o_2 _2867_ (.A1(\gen_pe[4].pe_inst.out_right[7] ),
    .A2(_0192_),
    .B1(_1543_),
    .B2(\gen_left[5][7] ),
    .C1(_2314_),
    .X(_0157_));
 sky130_fd_sc_hd__a22o_2 _2868_ (.A1(load),
    .A2(in_data_flat[168]),
    .B1(_0192_),
    .B2(\gen_pe[4].pe_inst.out_right[8] ),
    .X(_2315_));
 sky130_fd_sc_hd__a21o_2 _2869_ (.A1(\gen_left[5][8] ),
    .A2(_1543_),
    .B1(_2315_),
    .X(_0158_));
 sky130_fd_sc_hd__a22o_2 _2870_ (.A1(load),
    .A2(in_data_flat[169]),
    .B1(_0192_),
    .B2(\gen_pe[4].pe_inst.out_right[9] ),
    .X(_2316_));
 sky130_fd_sc_hd__a21o_2 _2871_ (.A1(\gen_left[5][9] ),
    .A2(_1543_),
    .B1(_2316_),
    .X(_0159_));
 sky130_fd_sc_hd__a22o_2 _2872_ (.A1(load),
    .A2(in_data_flat[170]),
    .B1(_0192_),
    .B2(\gen_pe[4].pe_inst.out_right[10] ),
    .X(_2317_));
 sky130_fd_sc_hd__a21o_2 _2873_ (.A1(\gen_left[5][10] ),
    .A2(_1543_),
    .B1(_2317_),
    .X(_0129_));
 sky130_fd_sc_hd__a22o_2 _2874_ (.A1(load),
    .A2(in_data_flat[171]),
    .B1(_0192_),
    .B2(\gen_pe[4].pe_inst.out_right[11] ),
    .X(_2318_));
 sky130_fd_sc_hd__a21o_2 _2875_ (.A1(\gen_left[5][11] ),
    .A2(_1543_),
    .B1(_2318_),
    .X(_0130_));
 sky130_fd_sc_hd__a22o_2 _2876_ (.A1(load),
    .A2(in_data_flat[172]),
    .B1(_0192_),
    .B2(\gen_pe[4].pe_inst.out_right[12] ),
    .X(_2319_));
 sky130_fd_sc_hd__a21o_2 _2877_ (.A1(\gen_left[5][12] ),
    .A2(_1543_),
    .B1(_2319_),
    .X(_0131_));
 sky130_fd_sc_hd__a22o_2 _2878_ (.A1(load),
    .A2(in_data_flat[173]),
    .B1(_0192_),
    .B2(\gen_pe[4].pe_inst.out_right[13] ),
    .X(_2320_));
 sky130_fd_sc_hd__a21o_2 _2879_ (.A1(\gen_left[5][13] ),
    .A2(_1543_),
    .B1(_2320_),
    .X(_0132_));
 sky130_fd_sc_hd__and2_2 _2880_ (.A(load),
    .B(in_data_flat[174]),
    .X(_2321_));
 sky130_fd_sc_hd__a221o_2 _2881_ (.A1(\gen_pe[4].pe_inst.out_right[14] ),
    .A2(_0192_),
    .B1(_1543_),
    .B2(\gen_left[5][14] ),
    .C1(_2321_),
    .X(_0133_));
 sky130_fd_sc_hd__and2_2 _2882_ (.A(load),
    .B(in_data_flat[175]),
    .X(_2322_));
 sky130_fd_sc_hd__a221o_2 _2883_ (.A1(\gen_pe[4].pe_inst.out_right[15] ),
    .A2(_0192_),
    .B1(_1543_),
    .B2(\gen_left[5][15] ),
    .C1(_2322_),
    .X(_0134_));
 sky130_fd_sc_hd__a22o_2 _2884_ (.A1(load),
    .A2(in_data_flat[176]),
    .B1(_0192_),
    .B2(\gen_pe[4].pe_inst.out_right[16] ),
    .X(_2323_));
 sky130_fd_sc_hd__a21o_2 _2885_ (.A1(\gen_left[5][16] ),
    .A2(_1543_),
    .B1(_2323_),
    .X(_0135_));
 sky130_fd_sc_hd__a22o_2 _2886_ (.A1(load),
    .A2(in_data_flat[177]),
    .B1(_0192_),
    .B2(\gen_pe[4].pe_inst.out_right[17] ),
    .X(_2324_));
 sky130_fd_sc_hd__a21o_2 _2887_ (.A1(\gen_left[5][17] ),
    .A2(_1543_),
    .B1(_2324_),
    .X(_0136_));
 sky130_fd_sc_hd__a22o_2 _2888_ (.A1(load),
    .A2(in_data_flat[178]),
    .B1(_0192_),
    .B2(\gen_pe[4].pe_inst.out_right[18] ),
    .X(_2325_));
 sky130_fd_sc_hd__a21o_2 _2889_ (.A1(\gen_left[5][18] ),
    .A2(_1543_),
    .B1(_2325_),
    .X(_0137_));
 sky130_fd_sc_hd__a22o_2 _2890_ (.A1(load),
    .A2(in_data_flat[179]),
    .B1(_0192_),
    .B2(\gen_pe[4].pe_inst.out_right[19] ),
    .X(_2326_));
 sky130_fd_sc_hd__a21o_2 _2891_ (.A1(\gen_left[5][19] ),
    .A2(_1543_),
    .B1(_2326_),
    .X(_0138_));
 sky130_fd_sc_hd__a22o_2 _2892_ (.A1(load),
    .A2(in_data_flat[180]),
    .B1(_0192_),
    .B2(\gen_pe[4].pe_inst.out_right[20] ),
    .X(_2327_));
 sky130_fd_sc_hd__a21o_2 _2893_ (.A1(\gen_left[5][20] ),
    .A2(_1543_),
    .B1(_2327_),
    .X(_0140_));
 sky130_fd_sc_hd__a22o_2 _2894_ (.A1(load),
    .A2(in_data_flat[181]),
    .B1(_0192_),
    .B2(\gen_pe[4].pe_inst.out_right[21] ),
    .X(_2328_));
 sky130_fd_sc_hd__a21o_2 _2895_ (.A1(\gen_left[5][21] ),
    .A2(_1543_),
    .B1(_2328_),
    .X(_0141_));
 sky130_fd_sc_hd__a22o_2 _2896_ (.A1(load),
    .A2(in_data_flat[182]),
    .B1(_0192_),
    .B2(\gen_pe[4].pe_inst.out_right[22] ),
    .X(_2329_));
 sky130_fd_sc_hd__a21o_2 _2897_ (.A1(\gen_left[5][22] ),
    .A2(_1543_),
    .B1(_2329_),
    .X(_0142_));
 sky130_fd_sc_hd__a22o_2 _2898_ (.A1(load),
    .A2(in_data_flat[183]),
    .B1(_0192_),
    .B2(\gen_pe[4].pe_inst.out_right[23] ),
    .X(_2330_));
 sky130_fd_sc_hd__a21o_2 _2899_ (.A1(\gen_left[5][23] ),
    .A2(_1543_),
    .B1(_2330_),
    .X(_0143_));
 sky130_fd_sc_hd__a22o_2 _2900_ (.A1(load),
    .A2(in_data_flat[184]),
    .B1(_0192_),
    .B2(\gen_pe[4].pe_inst.out_right[24] ),
    .X(_2331_));
 sky130_fd_sc_hd__a21o_2 _2901_ (.A1(\gen_left[5][24] ),
    .A2(_1543_),
    .B1(_2331_),
    .X(_0144_));
 sky130_fd_sc_hd__and2_2 _2902_ (.A(load),
    .B(in_data_flat[185]),
    .X(_2332_));
 sky130_fd_sc_hd__a221o_2 _2903_ (.A1(\gen_pe[4].pe_inst.out_right[25] ),
    .A2(_0192_),
    .B1(_1543_),
    .B2(\gen_left[5][25] ),
    .C1(_2332_),
    .X(_0145_));
 sky130_fd_sc_hd__a22o_2 _2904_ (.A1(load),
    .A2(in_data_flat[186]),
    .B1(_0192_),
    .B2(\gen_pe[4].pe_inst.out_right[26] ),
    .X(_2333_));
 sky130_fd_sc_hd__a21o_2 _2905_ (.A1(\gen_left[5][26] ),
    .A2(_1543_),
    .B1(_2333_),
    .X(_0146_));
 sky130_fd_sc_hd__a22o_2 _2906_ (.A1(load),
    .A2(in_data_flat[187]),
    .B1(_0192_),
    .B2(\gen_pe[4].pe_inst.out_right[27] ),
    .X(_2334_));
 sky130_fd_sc_hd__a21o_2 _2907_ (.A1(\gen_left[5][27] ),
    .A2(_1543_),
    .B1(_2334_),
    .X(_0147_));
 sky130_fd_sc_hd__and2_2 _2908_ (.A(load),
    .B(in_data_flat[188]),
    .X(_2335_));
 sky130_fd_sc_hd__a221o_2 _2909_ (.A1(\gen_pe[4].pe_inst.out_right[28] ),
    .A2(_0192_),
    .B1(_1543_),
    .B2(\gen_left[5][28] ),
    .C1(_2335_),
    .X(_0148_));
 sky130_fd_sc_hd__a22o_2 _2910_ (.A1(load),
    .A2(in_data_flat[189]),
    .B1(_0192_),
    .B2(\gen_pe[4].pe_inst.out_right[29] ),
    .X(_2336_));
 sky130_fd_sc_hd__a21o_2 _2911_ (.A1(\gen_left[5][29] ),
    .A2(_1543_),
    .B1(_2336_),
    .X(_0149_));
 sky130_fd_sc_hd__a22o_2 _2912_ (.A1(load),
    .A2(in_data_flat[190]),
    .B1(_0192_),
    .B2(\gen_pe[4].pe_inst.out_right[30] ),
    .X(_2337_));
 sky130_fd_sc_hd__a21o_2 _2913_ (.A1(\gen_left[5][30] ),
    .A2(_1543_),
    .B1(_2337_),
    .X(_0151_));
 sky130_fd_sc_hd__a22o_2 _2914_ (.A1(load),
    .A2(in_data_flat[191]),
    .B1(_0192_),
    .B2(\gen_pe[4].pe_inst.out_right[31] ),
    .X(_2338_));
 sky130_fd_sc_hd__a21o_2 _2915_ (.A1(\gen_left[5][31] ),
    .A2(_1543_),
    .B1(_2338_),
    .X(_0152_));
 sky130_fd_sc_hd__a22o_2 _2916_ (.A1(load),
    .A2(in_data_flat[192]),
    .B1(_0192_),
    .B2(\gen_left[6][0] ),
    .X(_2339_));
 sky130_fd_sc_hd__a21o_2 _2917_ (.A1(\gen_pe[5].pe_inst.out_right[0] ),
    .A2(_1543_),
    .B1(_2339_),
    .X(_0160_));
 sky130_fd_sc_hd__a22o_2 _2918_ (.A1(load),
    .A2(in_data_flat[193]),
    .B1(_0192_),
    .B2(\gen_left[6][1] ),
    .X(_2340_));
 sky130_fd_sc_hd__a21o_2 _2919_ (.A1(\gen_pe[5].pe_inst.out_right[1] ),
    .A2(_1543_),
    .B1(_2340_),
    .X(_0171_));
 sky130_fd_sc_hd__a22o_2 _2920_ (.A1(load),
    .A2(in_data_flat[194]),
    .B1(_0192_),
    .B2(\gen_left[6][2] ),
    .X(_2341_));
 sky130_fd_sc_hd__a21o_2 _2921_ (.A1(\gen_pe[5].pe_inst.out_right[2] ),
    .A2(_1543_),
    .B1(_2341_),
    .X(_0182_));
 sky130_fd_sc_hd__a22o_2 _2922_ (.A1(load),
    .A2(in_data_flat[195]),
    .B1(_0192_),
    .B2(\gen_left[6][3] ),
    .X(_2342_));
 sky130_fd_sc_hd__a21o_2 _2923_ (.A1(\gen_pe[5].pe_inst.out_right[3] ),
    .A2(_1543_),
    .B1(_2342_),
    .X(_0185_));
 sky130_fd_sc_hd__a22o_2 _2924_ (.A1(load),
    .A2(in_data_flat[196]),
    .B1(_0192_),
    .B2(\gen_left[6][4] ),
    .X(_2343_));
 sky130_fd_sc_hd__a21o_2 _2925_ (.A1(\gen_pe[5].pe_inst.out_right[4] ),
    .A2(_1543_),
    .B1(_2343_),
    .X(_0186_));
 sky130_fd_sc_hd__a22o_2 _2926_ (.A1(load),
    .A2(in_data_flat[197]),
    .B1(_0192_),
    .B2(\gen_left[6][5] ),
    .X(_2344_));
 sky130_fd_sc_hd__a21o_2 _2927_ (.A1(\gen_pe[5].pe_inst.out_right[5] ),
    .A2(_1543_),
    .B1(_2344_),
    .X(_0187_));
 sky130_fd_sc_hd__a22o_2 _2928_ (.A1(load),
    .A2(in_data_flat[198]),
    .B1(_0192_),
    .B2(\gen_left[6][6] ),
    .X(_2345_));
 sky130_fd_sc_hd__a21o_2 _2929_ (.A1(\gen_pe[5].pe_inst.out_right[6] ),
    .A2(_1543_),
    .B1(_2345_),
    .X(_0188_));
 sky130_fd_sc_hd__and2_2 _2930_ (.A(load),
    .B(in_data_flat[199]),
    .X(_2346_));
 sky130_fd_sc_hd__a221o_2 _2931_ (.A1(\gen_left[6][7] ),
    .A2(_0192_),
    .B1(_1543_),
    .B2(\gen_pe[5].pe_inst.out_right[7] ),
    .C1(_2346_),
    .X(_0189_));
 sky130_fd_sc_hd__a22o_2 _2932_ (.A1(load),
    .A2(in_data_flat[200]),
    .B1(_0192_),
    .B2(\gen_left[6][8] ),
    .X(_2347_));
 sky130_fd_sc_hd__a21o_2 _2933_ (.A1(\gen_pe[5].pe_inst.out_right[8] ),
    .A2(_1543_),
    .B1(_2347_),
    .X(_0190_));
 sky130_fd_sc_hd__a22o_2 _2934_ (.A1(load),
    .A2(in_data_flat[201]),
    .B1(_0192_),
    .B2(\gen_left[6][9] ),
    .X(_2348_));
 sky130_fd_sc_hd__a21o_2 _2935_ (.A1(\gen_pe[5].pe_inst.out_right[9] ),
    .A2(_1543_),
    .B1(_2348_),
    .X(_0191_));
 sky130_fd_sc_hd__a22o_2 _2936_ (.A1(load),
    .A2(in_data_flat[202]),
    .B1(_0192_),
    .B2(\gen_left[6][10] ),
    .X(_2349_));
 sky130_fd_sc_hd__a21o_2 _2937_ (.A1(\gen_pe[5].pe_inst.out_right[10] ),
    .A2(_1543_),
    .B1(_2349_),
    .X(_0161_));
 sky130_fd_sc_hd__a22o_2 _2938_ (.A1(load),
    .A2(in_data_flat[203]),
    .B1(_0192_),
    .B2(\gen_left[6][11] ),
    .X(_2350_));
 sky130_fd_sc_hd__a21o_2 _2939_ (.A1(\gen_pe[5].pe_inst.out_right[11] ),
    .A2(_1543_),
    .B1(_2350_),
    .X(_0162_));
 sky130_fd_sc_hd__a22o_2 _2940_ (.A1(load),
    .A2(in_data_flat[204]),
    .B1(_0192_),
    .B2(\gen_left[6][12] ),
    .X(_2351_));
 sky130_fd_sc_hd__a21o_2 _2941_ (.A1(\gen_pe[5].pe_inst.out_right[12] ),
    .A2(_1543_),
    .B1(_2351_),
    .X(_0163_));
 sky130_fd_sc_hd__a22o_2 _2942_ (.A1(load),
    .A2(in_data_flat[205]),
    .B1(_0192_),
    .B2(\gen_left[6][13] ),
    .X(_2352_));
 sky130_fd_sc_hd__a21o_2 _2943_ (.A1(\gen_pe[5].pe_inst.out_right[13] ),
    .A2(_1543_),
    .B1(_2352_),
    .X(_0164_));
 sky130_fd_sc_hd__and2_2 _2944_ (.A(load),
    .B(in_data_flat[206]),
    .X(_2353_));
 sky130_fd_sc_hd__a221o_2 _2945_ (.A1(\gen_left[6][14] ),
    .A2(_0192_),
    .B1(_1543_),
    .B2(\gen_pe[5].pe_inst.out_right[14] ),
    .C1(_2353_),
    .X(_0165_));
 sky130_fd_sc_hd__and2_2 _2946_ (.A(load),
    .B(in_data_flat[207]),
    .X(_2354_));
 sky130_fd_sc_hd__a221o_2 _2947_ (.A1(\gen_left[6][15] ),
    .A2(_0192_),
    .B1(_1543_),
    .B2(\gen_pe[5].pe_inst.out_right[15] ),
    .C1(_2354_),
    .X(_0166_));
 sky130_fd_sc_hd__a22o_2 _2948_ (.A1(load),
    .A2(in_data_flat[208]),
    .B1(_0192_),
    .B2(\gen_left[6][16] ),
    .X(_2355_));
 sky130_fd_sc_hd__a21o_2 _2949_ (.A1(\gen_pe[5].pe_inst.out_right[16] ),
    .A2(_1543_),
    .B1(_2355_),
    .X(_0167_));
 sky130_fd_sc_hd__a22o_2 _2950_ (.A1(load),
    .A2(in_data_flat[209]),
    .B1(_0192_),
    .B2(\gen_left[6][17] ),
    .X(_2356_));
 sky130_fd_sc_hd__a21o_2 _2951_ (.A1(\gen_pe[5].pe_inst.out_right[17] ),
    .A2(_1543_),
    .B1(_2356_),
    .X(_0168_));
 sky130_fd_sc_hd__a22o_2 _2952_ (.A1(load),
    .A2(in_data_flat[210]),
    .B1(_0192_),
    .B2(\gen_left[6][18] ),
    .X(_2357_));
 sky130_fd_sc_hd__a21o_2 _2953_ (.A1(\gen_pe[5].pe_inst.out_right[18] ),
    .A2(_1543_),
    .B1(_2357_),
    .X(_0169_));
 sky130_fd_sc_hd__a22o_2 _2954_ (.A1(load),
    .A2(in_data_flat[211]),
    .B1(_0192_),
    .B2(\gen_left[6][19] ),
    .X(_2358_));
 sky130_fd_sc_hd__a21o_2 _2955_ (.A1(\gen_pe[5].pe_inst.out_right[19] ),
    .A2(_1543_),
    .B1(_2358_),
    .X(_0170_));
 sky130_fd_sc_hd__a22o_2 _2956_ (.A1(load),
    .A2(in_data_flat[212]),
    .B1(_0192_),
    .B2(\gen_left[6][20] ),
    .X(_2359_));
 sky130_fd_sc_hd__a21o_2 _2957_ (.A1(\gen_pe[5].pe_inst.out_right[20] ),
    .A2(_1543_),
    .B1(_2359_),
    .X(_0172_));
 sky130_fd_sc_hd__a22o_2 _2958_ (.A1(load),
    .A2(in_data_flat[213]),
    .B1(_0192_),
    .B2(\gen_left[6][21] ),
    .X(_2360_));
 sky130_fd_sc_hd__a21o_2 _2959_ (.A1(\gen_pe[5].pe_inst.out_right[21] ),
    .A2(_1543_),
    .B1(_2360_),
    .X(_0173_));
 sky130_fd_sc_hd__a22o_2 _2960_ (.A1(load),
    .A2(in_data_flat[214]),
    .B1(_0192_),
    .B2(\gen_left[6][22] ),
    .X(_2361_));
 sky130_fd_sc_hd__a21o_2 _2961_ (.A1(\gen_pe[5].pe_inst.out_right[22] ),
    .A2(_1543_),
    .B1(_2361_),
    .X(_0174_));
 sky130_fd_sc_hd__a22o_2 _2962_ (.A1(load),
    .A2(in_data_flat[215]),
    .B1(_0192_),
    .B2(\gen_left[6][23] ),
    .X(_2362_));
 sky130_fd_sc_hd__a21o_2 _2963_ (.A1(\gen_pe[5].pe_inst.out_right[23] ),
    .A2(_1543_),
    .B1(_2362_),
    .X(_0175_));
 sky130_fd_sc_hd__a22o_2 _2964_ (.A1(load),
    .A2(in_data_flat[216]),
    .B1(_0192_),
    .B2(\gen_left[6][24] ),
    .X(_2363_));
 sky130_fd_sc_hd__a21o_2 _2965_ (.A1(\gen_pe[5].pe_inst.out_right[24] ),
    .A2(_1543_),
    .B1(_2363_),
    .X(_0176_));
 sky130_fd_sc_hd__and2_2 _2966_ (.A(load),
    .B(in_data_flat[217]),
    .X(_2364_));
 sky130_fd_sc_hd__a221o_2 _2967_ (.A1(\gen_left[6][25] ),
    .A2(_0192_),
    .B1(_1543_),
    .B2(\gen_pe[5].pe_inst.out_right[25] ),
    .C1(_2364_),
    .X(_0177_));
 sky130_fd_sc_hd__a22o_2 _2968_ (.A1(load),
    .A2(in_data_flat[218]),
    .B1(_0192_),
    .B2(\gen_left[6][26] ),
    .X(_2365_));
 sky130_fd_sc_hd__a21o_2 _2969_ (.A1(\gen_pe[5].pe_inst.out_right[26] ),
    .A2(_1543_),
    .B1(_2365_),
    .X(_0178_));
 sky130_fd_sc_hd__a22o_2 _2970_ (.A1(load),
    .A2(in_data_flat[219]),
    .B1(_0192_),
    .B2(\gen_left[6][27] ),
    .X(_2366_));
 sky130_fd_sc_hd__a21o_2 _2971_ (.A1(\gen_pe[5].pe_inst.out_right[27] ),
    .A2(_1543_),
    .B1(_2366_),
    .X(_0179_));
 sky130_fd_sc_hd__and2_2 _2972_ (.A(load),
    .B(in_data_flat[220]),
    .X(_2367_));
 sky130_fd_sc_hd__a221o_2 _2973_ (.A1(\gen_left[6][28] ),
    .A2(_0192_),
    .B1(_1543_),
    .B2(\gen_pe[5].pe_inst.out_right[28] ),
    .C1(_2367_),
    .X(_0180_));
 sky130_fd_sc_hd__a22o_2 _2974_ (.A1(load),
    .A2(in_data_flat[221]),
    .B1(_0192_),
    .B2(\gen_left[6][29] ),
    .X(_2368_));
 sky130_fd_sc_hd__a21o_2 _2975_ (.A1(\gen_pe[5].pe_inst.out_right[29] ),
    .A2(_1543_),
    .B1(_2368_),
    .X(_0181_));
 sky130_fd_sc_hd__a22o_2 _2976_ (.A1(load),
    .A2(in_data_flat[222]),
    .B1(_0192_),
    .B2(\gen_left[6][30] ),
    .X(_2369_));
 sky130_fd_sc_hd__a21o_2 _2977_ (.A1(\gen_pe[5].pe_inst.out_right[30] ),
    .A2(_1543_),
    .B1(_2369_),
    .X(_0183_));
 sky130_fd_sc_hd__a22o_2 _2978_ (.A1(load),
    .A2(in_data_flat[223]),
    .B1(_0192_),
    .B2(\gen_left[6][31] ),
    .X(_2370_));
 sky130_fd_sc_hd__a21o_2 _2979_ (.A1(\gen_pe[5].pe_inst.out_right[31] ),
    .A2(_1543_),
    .B1(_2370_),
    .X(_0184_));
 sky130_fd_sc_hd__inv_2 _2980_ (.A(rst),
    .Y(_0642_));
 sky130_fd_sc_hd__inv_2 _2981_ (.A(rst),
    .Y(_0643_));
 sky130_fd_sc_hd__inv_2 _2982_ (.A(rst),
    .Y(_0644_));
 sky130_fd_sc_hd__inv_2 _2983_ (.A(rst),
    .Y(_0645_));
 sky130_fd_sc_hd__inv_2 _2984_ (.A(rst),
    .Y(_0646_));
 sky130_fd_sc_hd__inv_2 _2985_ (.A(rst),
    .Y(_0647_));
 sky130_fd_sc_hd__inv_2 _2986_ (.A(rst),
    .Y(_0648_));
 sky130_fd_sc_hd__inv_2 _2987_ (.A(rst),
    .Y(_0649_));
 sky130_fd_sc_hd__inv_2 _2988_ (.A(rst),
    .Y(_0650_));
 sky130_fd_sc_hd__inv_2 _2989_ (.A(rst),
    .Y(_0651_));
 sky130_fd_sc_hd__inv_2 _2990_ (.A(rst),
    .Y(_0652_));
 sky130_fd_sc_hd__inv_2 _2991_ (.A(rst),
    .Y(_0653_));
 sky130_fd_sc_hd__inv_2 _2992_ (.A(rst),
    .Y(_0654_));
 sky130_fd_sc_hd__inv_2 _2993_ (.A(rst),
    .Y(_0655_));
 sky130_fd_sc_hd__inv_2 _2994_ (.A(rst),
    .Y(_0656_));
 sky130_fd_sc_hd__inv_2 _2995_ (.A(rst),
    .Y(_0657_));
 sky130_fd_sc_hd__inv_2 _2996_ (.A(rst),
    .Y(_0658_));
 sky130_fd_sc_hd__inv_2 _2997_ (.A(rst),
    .Y(_0659_));
 sky130_fd_sc_hd__inv_2 _2998_ (.A(rst),
    .Y(_0660_));
 sky130_fd_sc_hd__inv_2 _2999_ (.A(rst),
    .Y(_0661_));
 sky130_fd_sc_hd__inv_2 _3000_ (.A(rst),
    .Y(_0662_));
 sky130_fd_sc_hd__inv_2 _3001_ (.A(rst),
    .Y(_0663_));
 sky130_fd_sc_hd__inv_2 _3002_ (.A(rst),
    .Y(_0664_));
 sky130_fd_sc_hd__inv_2 _3003_ (.A(rst),
    .Y(_0665_));
 sky130_fd_sc_hd__inv_2 _3004_ (.A(rst),
    .Y(_0666_));
 sky130_fd_sc_hd__inv_2 _3005_ (.A(rst),
    .Y(_0667_));
 sky130_fd_sc_hd__inv_2 _3006_ (.A(rst),
    .Y(_0668_));
 sky130_fd_sc_hd__inv_2 _3007_ (.A(rst),
    .Y(_0669_));
 sky130_fd_sc_hd__inv_2 _3008_ (.A(rst),
    .Y(_0670_));
 sky130_fd_sc_hd__inv_2 _3009_ (.A(rst),
    .Y(_0671_));
 sky130_fd_sc_hd__inv_2 _3010_ (.A(rst),
    .Y(_0672_));
 sky130_fd_sc_hd__inv_2 _3011_ (.A(rst),
    .Y(_0673_));
 sky130_fd_sc_hd__inv_2 _3012_ (.A(rst),
    .Y(_0674_));
 sky130_fd_sc_hd__inv_2 _3013_ (.A(rst),
    .Y(_0675_));
 sky130_fd_sc_hd__inv_2 _3014_ (.A(rst),
    .Y(_0676_));
 sky130_fd_sc_hd__inv_2 _3015_ (.A(rst),
    .Y(_0677_));
 sky130_fd_sc_hd__inv_2 _3016_ (.A(rst),
    .Y(_0678_));
 sky130_fd_sc_hd__inv_2 _3017_ (.A(rst),
    .Y(_0679_));
 sky130_fd_sc_hd__inv_2 _3018_ (.A(rst),
    .Y(_0680_));
 sky130_fd_sc_hd__inv_2 _3019_ (.A(rst),
    .Y(_0681_));
 sky130_fd_sc_hd__inv_2 _3020_ (.A(rst),
    .Y(_0682_));
 sky130_fd_sc_hd__inv_2 _3021_ (.A(rst),
    .Y(_0683_));
 sky130_fd_sc_hd__inv_2 _3022_ (.A(rst),
    .Y(_0684_));
 sky130_fd_sc_hd__inv_2 _3023_ (.A(rst),
    .Y(_0685_));
 sky130_fd_sc_hd__inv_2 _3024_ (.A(rst),
    .Y(_0686_));
 sky130_fd_sc_hd__inv_2 _3025_ (.A(rst),
    .Y(_0687_));
 sky130_fd_sc_hd__inv_2 _3026_ (.A(rst),
    .Y(_0688_));
 sky130_fd_sc_hd__inv_2 _3027_ (.A(rst),
    .Y(_0689_));
 sky130_fd_sc_hd__inv_2 _3028_ (.A(rst),
    .Y(_0690_));
 sky130_fd_sc_hd__inv_2 _3029_ (.A(rst),
    .Y(_0691_));
 sky130_fd_sc_hd__inv_2 _3030_ (.A(rst),
    .Y(_0692_));
 sky130_fd_sc_hd__inv_2 _3031_ (.A(rst),
    .Y(_0693_));
 sky130_fd_sc_hd__inv_2 _3032_ (.A(rst),
    .Y(_0694_));
 sky130_fd_sc_hd__inv_2 _3033_ (.A(rst),
    .Y(_0695_));
 sky130_fd_sc_hd__inv_2 _3034_ (.A(rst),
    .Y(_0696_));
 sky130_fd_sc_hd__inv_2 _3035_ (.A(rst),
    .Y(_0697_));
 sky130_fd_sc_hd__inv_2 _3036_ (.A(rst),
    .Y(_0698_));
 sky130_fd_sc_hd__inv_2 _3037_ (.A(rst),
    .Y(_0699_));
 sky130_fd_sc_hd__inv_2 _3038_ (.A(rst),
    .Y(_0700_));
 sky130_fd_sc_hd__inv_2 _3039_ (.A(rst),
    .Y(_0701_));
 sky130_fd_sc_hd__inv_2 _3040_ (.A(rst),
    .Y(_0702_));
 sky130_fd_sc_hd__inv_2 _3041_ (.A(rst),
    .Y(_0703_));
 sky130_fd_sc_hd__inv_2 _3042_ (.A(rst),
    .Y(_0704_));
 sky130_fd_sc_hd__inv_2 _3043_ (.A(rst),
    .Y(_0705_));
 sky130_fd_sc_hd__inv_2 _3044_ (.A(rst),
    .Y(_0706_));
 sky130_fd_sc_hd__inv_2 _3045_ (.A(rst),
    .Y(_0707_));
 sky130_fd_sc_hd__inv_2 _3046_ (.A(rst),
    .Y(_0708_));
 sky130_fd_sc_hd__inv_2 _3047_ (.A(rst),
    .Y(_0709_));
 sky130_fd_sc_hd__inv_2 _3048_ (.A(rst),
    .Y(_0710_));
 sky130_fd_sc_hd__inv_2 _3049_ (.A(rst),
    .Y(_0711_));
 sky130_fd_sc_hd__inv_2 _3050_ (.A(rst),
    .Y(_0712_));
 sky130_fd_sc_hd__inv_2 _3051_ (.A(rst),
    .Y(_0713_));
 sky130_fd_sc_hd__inv_2 _3052_ (.A(rst),
    .Y(_0714_));
 sky130_fd_sc_hd__inv_2 _3053_ (.A(rst),
    .Y(_0715_));
 sky130_fd_sc_hd__inv_2 _3054_ (.A(rst),
    .Y(_0716_));
 sky130_fd_sc_hd__inv_2 _3055_ (.A(rst),
    .Y(_0717_));
 sky130_fd_sc_hd__inv_2 _3056_ (.A(rst),
    .Y(_0718_));
 sky130_fd_sc_hd__inv_2 _3057_ (.A(rst),
    .Y(_0719_));
 sky130_fd_sc_hd__inv_2 _3058_ (.A(rst),
    .Y(_0720_));
 sky130_fd_sc_hd__inv_2 _3059_ (.A(rst),
    .Y(_0721_));
 sky130_fd_sc_hd__inv_2 _3060_ (.A(rst),
    .Y(_0722_));
 sky130_fd_sc_hd__inv_2 _3061_ (.A(rst),
    .Y(_0723_));
 sky130_fd_sc_hd__inv_2 _3062_ (.A(rst),
    .Y(_0724_));
 sky130_fd_sc_hd__inv_2 _3063_ (.A(rst),
    .Y(_0725_));
 sky130_fd_sc_hd__inv_2 _3064_ (.A(rst),
    .Y(_0726_));
 sky130_fd_sc_hd__inv_2 _3065_ (.A(rst),
    .Y(_0727_));
 sky130_fd_sc_hd__inv_2 _3066_ (.A(rst),
    .Y(_0728_));
 sky130_fd_sc_hd__inv_2 _3067_ (.A(rst),
    .Y(_0729_));
 sky130_fd_sc_hd__inv_2 _3068_ (.A(rst),
    .Y(_0730_));
 sky130_fd_sc_hd__inv_2 _3069_ (.A(rst),
    .Y(_0731_));
 sky130_fd_sc_hd__inv_2 _3070_ (.A(rst),
    .Y(_0732_));
 sky130_fd_sc_hd__inv_2 _3071_ (.A(rst),
    .Y(_0733_));
 sky130_fd_sc_hd__inv_2 _3072_ (.A(rst),
    .Y(_0734_));
 sky130_fd_sc_hd__inv_2 _3073_ (.A(rst),
    .Y(_0735_));
 sky130_fd_sc_hd__inv_2 _3074_ (.A(rst),
    .Y(_0736_));
 sky130_fd_sc_hd__inv_2 _3075_ (.A(rst),
    .Y(_0737_));
 sky130_fd_sc_hd__inv_2 _3076_ (.A(rst),
    .Y(_0738_));
 sky130_fd_sc_hd__inv_2 _3077_ (.A(rst),
    .Y(_0739_));
 sky130_fd_sc_hd__inv_2 _3078_ (.A(rst),
    .Y(_0740_));
 sky130_fd_sc_hd__inv_2 _3079_ (.A(rst),
    .Y(_0741_));
 sky130_fd_sc_hd__inv_2 _3080_ (.A(rst),
    .Y(_0742_));
 sky130_fd_sc_hd__inv_2 _3081_ (.A(rst),
    .Y(_0743_));
 sky130_fd_sc_hd__inv_2 _3082_ (.A(rst),
    .Y(_0744_));
 sky130_fd_sc_hd__inv_2 _3083_ (.A(rst),
    .Y(_0745_));
 sky130_fd_sc_hd__inv_2 _3084_ (.A(rst),
    .Y(_0746_));
 sky130_fd_sc_hd__inv_2 _3085_ (.A(rst),
    .Y(_0747_));
 sky130_fd_sc_hd__inv_2 _3086_ (.A(rst),
    .Y(_0748_));
 sky130_fd_sc_hd__inv_2 _3087_ (.A(rst),
    .Y(_0749_));
 sky130_fd_sc_hd__inv_2 _3088_ (.A(rst),
    .Y(_0750_));
 sky130_fd_sc_hd__inv_2 _3089_ (.A(rst),
    .Y(_0751_));
 sky130_fd_sc_hd__inv_2 _3090_ (.A(rst),
    .Y(_0752_));
 sky130_fd_sc_hd__inv_2 _3091_ (.A(rst),
    .Y(_0753_));
 sky130_fd_sc_hd__inv_2 _3092_ (.A(rst),
    .Y(_0754_));
 sky130_fd_sc_hd__inv_2 _3093_ (.A(rst),
    .Y(_0755_));
 sky130_fd_sc_hd__inv_2 _3094_ (.A(rst),
    .Y(_0756_));
 sky130_fd_sc_hd__inv_2 _3095_ (.A(rst),
    .Y(_0757_));
 sky130_fd_sc_hd__inv_2 _3096_ (.A(rst),
    .Y(_0758_));
 sky130_fd_sc_hd__inv_2 _3097_ (.A(rst),
    .Y(_0759_));
 sky130_fd_sc_hd__inv_2 _3098_ (.A(rst),
    .Y(_0760_));
 sky130_fd_sc_hd__inv_2 _3099_ (.A(rst),
    .Y(_0761_));
 sky130_fd_sc_hd__inv_2 _3100_ (.A(rst),
    .Y(_0762_));
 sky130_fd_sc_hd__inv_2 _3101_ (.A(rst),
    .Y(_0763_));
 sky130_fd_sc_hd__inv_2 _3102_ (.A(rst),
    .Y(_0764_));
 sky130_fd_sc_hd__inv_2 _3103_ (.A(rst),
    .Y(_0765_));
 sky130_fd_sc_hd__inv_2 _3104_ (.A(rst),
    .Y(_0766_));
 sky130_fd_sc_hd__inv_2 _3105_ (.A(rst),
    .Y(_0767_));
 sky130_fd_sc_hd__inv_2 _3106_ (.A(rst),
    .Y(_0768_));
 sky130_fd_sc_hd__inv_2 _3107_ (.A(rst),
    .Y(_0769_));
 sky130_fd_sc_hd__inv_2 _3108_ (.A(rst),
    .Y(_0770_));
 sky130_fd_sc_hd__inv_2 _3109_ (.A(rst),
    .Y(_0771_));
 sky130_fd_sc_hd__inv_2 _3110_ (.A(rst),
    .Y(_0772_));
 sky130_fd_sc_hd__inv_2 _3111_ (.A(rst),
    .Y(_0773_));
 sky130_fd_sc_hd__inv_2 _3112_ (.A(rst),
    .Y(_0774_));
 sky130_fd_sc_hd__inv_2 _3113_ (.A(rst),
    .Y(_0775_));
 sky130_fd_sc_hd__inv_2 _3114_ (.A(rst),
    .Y(_0776_));
 sky130_fd_sc_hd__inv_2 _3115_ (.A(rst),
    .Y(_0777_));
 sky130_fd_sc_hd__inv_2 _3116_ (.A(rst),
    .Y(_0778_));
 sky130_fd_sc_hd__inv_2 _3117_ (.A(rst),
    .Y(_0779_));
 sky130_fd_sc_hd__inv_2 _3118_ (.A(rst),
    .Y(_0780_));
 sky130_fd_sc_hd__inv_2 _3119_ (.A(rst),
    .Y(_0781_));
 sky130_fd_sc_hd__inv_2 _3120_ (.A(rst),
    .Y(_0782_));
 sky130_fd_sc_hd__inv_2 _3121_ (.A(rst),
    .Y(_0783_));
 sky130_fd_sc_hd__inv_2 _3122_ (.A(rst),
    .Y(_0784_));
 sky130_fd_sc_hd__inv_2 _3123_ (.A(rst),
    .Y(_0785_));
 sky130_fd_sc_hd__inv_2 _3124_ (.A(rst),
    .Y(_0786_));
 sky130_fd_sc_hd__inv_2 _3125_ (.A(rst),
    .Y(_0787_));
 sky130_fd_sc_hd__inv_2 _3126_ (.A(rst),
    .Y(_0788_));
 sky130_fd_sc_hd__inv_2 _3127_ (.A(rst),
    .Y(_0789_));
 sky130_fd_sc_hd__inv_2 _3128_ (.A(rst),
    .Y(_0790_));
 sky130_fd_sc_hd__inv_2 _3129_ (.A(rst),
    .Y(_0791_));
 sky130_fd_sc_hd__inv_2 _3130_ (.A(rst),
    .Y(_0792_));
 sky130_fd_sc_hd__inv_2 _3131_ (.A(rst),
    .Y(_0793_));
 sky130_fd_sc_hd__inv_2 _3132_ (.A(rst),
    .Y(_0794_));
 sky130_fd_sc_hd__inv_2 _3133_ (.A(rst),
    .Y(_0795_));
 sky130_fd_sc_hd__inv_2 _3134_ (.A(rst),
    .Y(_0796_));
 sky130_fd_sc_hd__inv_2 _3135_ (.A(rst),
    .Y(_0797_));
 sky130_fd_sc_hd__inv_2 _3136_ (.A(rst),
    .Y(_0798_));
 sky130_fd_sc_hd__inv_2 _3137_ (.A(rst),
    .Y(_0799_));
 sky130_fd_sc_hd__inv_2 _3138_ (.A(rst),
    .Y(_0800_));
 sky130_fd_sc_hd__inv_2 _3139_ (.A(rst),
    .Y(_0801_));
 sky130_fd_sc_hd__inv_2 _3140_ (.A(rst),
    .Y(_0802_));
 sky130_fd_sc_hd__inv_2 _3141_ (.A(rst),
    .Y(_0803_));
 sky130_fd_sc_hd__inv_2 _3142_ (.A(rst),
    .Y(_0804_));
 sky130_fd_sc_hd__inv_2 _3143_ (.A(rst),
    .Y(_0805_));
 sky130_fd_sc_hd__inv_2 _3144_ (.A(rst),
    .Y(_0806_));
 sky130_fd_sc_hd__inv_2 _3145_ (.A(rst),
    .Y(_0807_));
 sky130_fd_sc_hd__inv_2 _3146_ (.A(rst),
    .Y(_0808_));
 sky130_fd_sc_hd__inv_2 _3147_ (.A(rst),
    .Y(_0809_));
 sky130_fd_sc_hd__inv_2 _3148_ (.A(rst),
    .Y(_0810_));
 sky130_fd_sc_hd__inv_2 _3149_ (.A(rst),
    .Y(_0811_));
 sky130_fd_sc_hd__inv_2 _3150_ (.A(rst),
    .Y(_0812_));
 sky130_fd_sc_hd__inv_2 _3151_ (.A(rst),
    .Y(_0813_));
 sky130_fd_sc_hd__inv_2 _3152_ (.A(rst),
    .Y(_0814_));
 sky130_fd_sc_hd__inv_2 _3153_ (.A(rst),
    .Y(_0815_));
 sky130_fd_sc_hd__inv_2 _3154_ (.A(rst),
    .Y(_0816_));
 sky130_fd_sc_hd__inv_2 _3155_ (.A(rst),
    .Y(_0817_));
 sky130_fd_sc_hd__inv_2 _3156_ (.A(rst),
    .Y(_0818_));
 sky130_fd_sc_hd__inv_2 _3157_ (.A(rst),
    .Y(_0819_));
 sky130_fd_sc_hd__inv_2 _3158_ (.A(rst),
    .Y(_0820_));
 sky130_fd_sc_hd__inv_2 _3159_ (.A(rst),
    .Y(_0821_));
 sky130_fd_sc_hd__inv_2 _3160_ (.A(rst),
    .Y(_0822_));
 sky130_fd_sc_hd__inv_2 _3161_ (.A(rst),
    .Y(_0823_));
 sky130_fd_sc_hd__inv_2 _3162_ (.A(rst),
    .Y(_0824_));
 sky130_fd_sc_hd__inv_2 _3163_ (.A(rst),
    .Y(_0825_));
 sky130_fd_sc_hd__inv_2 _3164_ (.A(rst),
    .Y(_0826_));
 sky130_fd_sc_hd__inv_2 _3165_ (.A(rst),
    .Y(_0827_));
 sky130_fd_sc_hd__inv_2 _3166_ (.A(rst),
    .Y(_0828_));
 sky130_fd_sc_hd__inv_2 _3167_ (.A(rst),
    .Y(_0829_));
 sky130_fd_sc_hd__inv_2 _3168_ (.A(rst),
    .Y(_0830_));
 sky130_fd_sc_hd__inv_2 _3169_ (.A(rst),
    .Y(_0831_));
 sky130_fd_sc_hd__inv_2 _3170_ (.A(rst),
    .Y(_0832_));
 sky130_fd_sc_hd__inv_2 _3171_ (.A(rst),
    .Y(_0833_));
 sky130_fd_sc_hd__inv_2 _3172_ (.A(rst),
    .Y(_0834_));
 sky130_fd_sc_hd__inv_2 _3173_ (.A(rst),
    .Y(_0835_));
 sky130_fd_sc_hd__inv_2 _3174_ (.A(rst),
    .Y(_0836_));
 sky130_fd_sc_hd__inv_2 _3175_ (.A(rst),
    .Y(_0837_));
 sky130_fd_sc_hd__inv_2 _3176_ (.A(rst),
    .Y(_0838_));
 sky130_fd_sc_hd__inv_2 _3177_ (.A(rst),
    .Y(_0839_));
 sky130_fd_sc_hd__inv_2 _3178_ (.A(rst),
    .Y(_0840_));
 sky130_fd_sc_hd__inv_2 _3179_ (.A(rst),
    .Y(_0841_));
 sky130_fd_sc_hd__inv_2 _3180_ (.A(rst),
    .Y(_0842_));
 sky130_fd_sc_hd__inv_2 _3181_ (.A(rst),
    .Y(_0843_));
 sky130_fd_sc_hd__inv_2 _3182_ (.A(rst),
    .Y(_0844_));
 sky130_fd_sc_hd__inv_2 _3183_ (.A(rst),
    .Y(_0845_));
 sky130_fd_sc_hd__inv_2 _3184_ (.A(rst),
    .Y(_0846_));
 sky130_fd_sc_hd__inv_2 _3185_ (.A(rst),
    .Y(_0847_));
 sky130_fd_sc_hd__inv_2 _3186_ (.A(rst),
    .Y(_0848_));
 sky130_fd_sc_hd__inv_2 _3187_ (.A(rst),
    .Y(_0849_));
 sky130_fd_sc_hd__inv_2 _3188_ (.A(rst),
    .Y(_0850_));
 sky130_fd_sc_hd__inv_2 _3189_ (.A(rst),
    .Y(_0851_));
 sky130_fd_sc_hd__inv_2 _3190_ (.A(rst),
    .Y(_0852_));
 sky130_fd_sc_hd__inv_2 _3191_ (.A(rst),
    .Y(_0853_));
 sky130_fd_sc_hd__inv_2 _3192_ (.A(rst),
    .Y(_0854_));
 sky130_fd_sc_hd__inv_2 _3193_ (.A(rst),
    .Y(_0855_));
 sky130_fd_sc_hd__inv_2 _3194_ (.A(rst),
    .Y(_0856_));
 sky130_fd_sc_hd__inv_2 _3195_ (.A(rst),
    .Y(_0857_));
 sky130_fd_sc_hd__inv_2 _3196_ (.A(rst),
    .Y(_0858_));
 sky130_fd_sc_hd__inv_2 _3197_ (.A(rst),
    .Y(_0859_));
 sky130_fd_sc_hd__inv_2 _3198_ (.A(rst),
    .Y(_0860_));
 sky130_fd_sc_hd__inv_2 _3199_ (.A(rst),
    .Y(_0861_));
 sky130_fd_sc_hd__inv_2 _3200_ (.A(rst),
    .Y(_0862_));
 sky130_fd_sc_hd__inv_2 _3201_ (.A(rst),
    .Y(_0863_));
 sky130_fd_sc_hd__inv_2 _3202_ (.A(rst),
    .Y(_0864_));
 sky130_fd_sc_hd__inv_2 _3203_ (.A(rst),
    .Y(_0865_));
 sky130_fd_sc_hd__inv_2 _3204_ (.A(rst),
    .Y(_0866_));
 sky130_fd_sc_hd__inv_2 _3205_ (.A(rst),
    .Y(_0867_));
 sky130_fd_sc_hd__inv_2 _3206_ (.A(rst),
    .Y(_0868_));
 sky130_fd_sc_hd__inv_2 _3207_ (.A(rst),
    .Y(_0869_));
 sky130_fd_sc_hd__inv_2 _3208_ (.A(rst),
    .Y(_0870_));
 sky130_fd_sc_hd__inv_2 _3209_ (.A(rst),
    .Y(_0871_));
 sky130_fd_sc_hd__inv_2 _3210_ (.A(rst),
    .Y(_0872_));
 sky130_fd_sc_hd__inv_2 _3211_ (.A(rst),
    .Y(_0873_));
 sky130_fd_sc_hd__inv_2 _3212_ (.A(rst),
    .Y(_0874_));
 sky130_fd_sc_hd__inv_2 _3213_ (.A(rst),
    .Y(_0875_));
 sky130_fd_sc_hd__inv_2 _3214_ (.A(rst),
    .Y(_0876_));
 sky130_fd_sc_hd__inv_2 _3215_ (.A(rst),
    .Y(_0877_));
 sky130_fd_sc_hd__inv_2 _3216_ (.A(rst),
    .Y(_0878_));
 sky130_fd_sc_hd__inv_2 _3217_ (.A(rst),
    .Y(_0879_));
 sky130_fd_sc_hd__inv_2 _3218_ (.A(rst),
    .Y(_0880_));
 sky130_fd_sc_hd__inv_2 _3219_ (.A(rst),
    .Y(_0881_));
 sky130_fd_sc_hd__inv_2 _3220_ (.A(rst),
    .Y(_0882_));
 sky130_fd_sc_hd__inv_2 _3221_ (.A(rst),
    .Y(_0883_));
 sky130_fd_sc_hd__inv_2 _3222_ (.A(rst),
    .Y(_0884_));
 sky130_fd_sc_hd__inv_2 _3223_ (.A(rst),
    .Y(_0885_));
 sky130_fd_sc_hd__inv_2 _3224_ (.A(rst),
    .Y(_0886_));
 sky130_fd_sc_hd__inv_2 _3225_ (.A(rst),
    .Y(_0887_));
 sky130_fd_sc_hd__inv_2 _3226_ (.A(rst),
    .Y(_0888_));
 sky130_fd_sc_hd__inv_2 _3227_ (.A(rst),
    .Y(_0889_));
 sky130_fd_sc_hd__inv_2 _3228_ (.A(rst),
    .Y(_0890_));
 sky130_fd_sc_hd__inv_2 _3229_ (.A(rst),
    .Y(_0891_));
 sky130_fd_sc_hd__inv_2 _3230_ (.A(rst),
    .Y(_0892_));
 sky130_fd_sc_hd__inv_2 _3231_ (.A(rst),
    .Y(_0893_));
 sky130_fd_sc_hd__inv_2 _3232_ (.A(rst),
    .Y(_0894_));
 sky130_fd_sc_hd__inv_2 _3233_ (.A(rst),
    .Y(_0895_));
 sky130_fd_sc_hd__inv_2 _3234_ (.A(rst),
    .Y(_0896_));
 sky130_fd_sc_hd__inv_2 _3235_ (.A(rst),
    .Y(_0897_));
 sky130_fd_sc_hd__inv_2 _3236_ (.A(rst),
    .Y(_0898_));
 sky130_fd_sc_hd__inv_2 _3237_ (.A(rst),
    .Y(_0899_));
 sky130_fd_sc_hd__inv_2 _3238_ (.A(rst),
    .Y(_0900_));
 sky130_fd_sc_hd__inv_2 _3239_ (.A(rst),
    .Y(_0901_));
 sky130_fd_sc_hd__inv_2 _3240_ (.A(rst),
    .Y(_0902_));
 sky130_fd_sc_hd__inv_2 _3241_ (.A(rst),
    .Y(_0903_));
 sky130_fd_sc_hd__inv_2 _3242_ (.A(rst),
    .Y(_0904_));
 sky130_fd_sc_hd__inv_2 _3243_ (.A(rst),
    .Y(_0905_));
 sky130_fd_sc_hd__inv_2 _3244_ (.A(rst),
    .Y(_0906_));
 sky130_fd_sc_hd__inv_2 _3245_ (.A(rst),
    .Y(_0907_));
 sky130_fd_sc_hd__inv_2 _3246_ (.A(rst),
    .Y(_0908_));
 sky130_fd_sc_hd__inv_2 _3247_ (.A(rst),
    .Y(_0909_));
 sky130_fd_sc_hd__inv_2 _3248_ (.A(rst),
    .Y(_0910_));
 sky130_fd_sc_hd__inv_2 _3249_ (.A(rst),
    .Y(_0911_));
 sky130_fd_sc_hd__inv_2 _3250_ (.A(rst),
    .Y(_0912_));
 sky130_fd_sc_hd__inv_2 _3251_ (.A(rst),
    .Y(_0913_));
 sky130_fd_sc_hd__inv_2 _3252_ (.A(rst),
    .Y(_0914_));
 sky130_fd_sc_hd__inv_2 _3253_ (.A(rst),
    .Y(_0915_));
 sky130_fd_sc_hd__inv_2 _3254_ (.A(rst),
    .Y(_0916_));
 sky130_fd_sc_hd__inv_2 _3255_ (.A(rst),
    .Y(_0917_));
 sky130_fd_sc_hd__inv_2 _3256_ (.A(rst),
    .Y(_0918_));
 sky130_fd_sc_hd__inv_2 _3257_ (.A(rst),
    .Y(_0919_));
 sky130_fd_sc_hd__inv_2 _3258_ (.A(rst),
    .Y(_0920_));
 sky130_fd_sc_hd__inv_2 _3259_ (.A(rst),
    .Y(_0921_));
 sky130_fd_sc_hd__inv_2 _3260_ (.A(rst),
    .Y(_0922_));
 sky130_fd_sc_hd__inv_2 _3261_ (.A(rst),
    .Y(_0923_));
 sky130_fd_sc_hd__inv_2 _3262_ (.A(rst),
    .Y(_0924_));
 sky130_fd_sc_hd__inv_2 _3263_ (.A(rst),
    .Y(_0925_));
 sky130_fd_sc_hd__inv_2 _3264_ (.A(rst),
    .Y(_0926_));
 sky130_fd_sc_hd__inv_2 _3265_ (.A(rst),
    .Y(_0927_));
 sky130_fd_sc_hd__inv_2 _3266_ (.A(rst),
    .Y(_0928_));
 sky130_fd_sc_hd__inv_2 _3267_ (.A(rst),
    .Y(_0929_));
 sky130_fd_sc_hd__inv_2 _3268_ (.A(rst),
    .Y(_0930_));
 sky130_fd_sc_hd__inv_2 _3269_ (.A(rst),
    .Y(_0931_));
 sky130_fd_sc_hd__inv_2 _3270_ (.A(rst),
    .Y(_0932_));
 sky130_fd_sc_hd__inv_2 _3271_ (.A(rst),
    .Y(_0933_));
 sky130_fd_sc_hd__inv_2 _3272_ (.A(rst),
    .Y(_0934_));
 sky130_fd_sc_hd__inv_2 _3273_ (.A(rst),
    .Y(_0935_));
 sky130_fd_sc_hd__inv_2 _3274_ (.A(rst),
    .Y(_0936_));
 sky130_fd_sc_hd__inv_2 _3275_ (.A(rst),
    .Y(_0937_));
 sky130_fd_sc_hd__inv_2 _3276_ (.A(rst),
    .Y(_0938_));
 sky130_fd_sc_hd__inv_2 _3277_ (.A(rst),
    .Y(_0939_));
 sky130_fd_sc_hd__inv_2 _3278_ (.A(rst),
    .Y(_0940_));
 sky130_fd_sc_hd__inv_2 _3279_ (.A(rst),
    .Y(_0941_));
 sky130_fd_sc_hd__inv_2 _3280_ (.A(rst),
    .Y(_0942_));
 sky130_fd_sc_hd__inv_2 _3281_ (.A(rst),
    .Y(_0943_));
 sky130_fd_sc_hd__inv_2 _3282_ (.A(rst),
    .Y(_0944_));
 sky130_fd_sc_hd__inv_2 _3283_ (.A(rst),
    .Y(_0945_));
 sky130_fd_sc_hd__inv_2 _3284_ (.A(rst),
    .Y(_0946_));
 sky130_fd_sc_hd__inv_2 _3285_ (.A(rst),
    .Y(_0947_));
 sky130_fd_sc_hd__inv_2 _3286_ (.A(rst),
    .Y(_0948_));
 sky130_fd_sc_hd__inv_2 _3287_ (.A(rst),
    .Y(_0949_));
 sky130_fd_sc_hd__inv_2 _3288_ (.A(rst),
    .Y(_0950_));
 sky130_fd_sc_hd__inv_2 _3289_ (.A(rst),
    .Y(_0951_));
 sky130_fd_sc_hd__inv_2 _3290_ (.A(rst),
    .Y(_0952_));
 sky130_fd_sc_hd__inv_2 _3291_ (.A(rst),
    .Y(_0953_));
 sky130_fd_sc_hd__inv_2 _3292_ (.A(rst),
    .Y(_0954_));
 sky130_fd_sc_hd__inv_2 _3293_ (.A(rst),
    .Y(_0955_));
 sky130_fd_sc_hd__inv_2 _3294_ (.A(rst),
    .Y(_0956_));
 sky130_fd_sc_hd__inv_2 _3295_ (.A(rst),
    .Y(_0957_));
 sky130_fd_sc_hd__inv_2 _3296_ (.A(rst),
    .Y(_0958_));
 sky130_fd_sc_hd__inv_2 _3297_ (.A(rst),
    .Y(_0959_));
 sky130_fd_sc_hd__inv_2 _3298_ (.A(rst),
    .Y(_0960_));
 sky130_fd_sc_hd__inv_2 _3299_ (.A(rst),
    .Y(_0961_));
 sky130_fd_sc_hd__inv_2 _3300_ (.A(rst),
    .Y(_0962_));
 sky130_fd_sc_hd__inv_2 _3301_ (.A(rst),
    .Y(_0963_));
 sky130_fd_sc_hd__inv_2 _3302_ (.A(rst),
    .Y(_0964_));
 sky130_fd_sc_hd__inv_2 _3303_ (.A(rst),
    .Y(_0965_));
 sky130_fd_sc_hd__inv_2 _3304_ (.A(rst),
    .Y(_0966_));
 sky130_fd_sc_hd__inv_2 _3305_ (.A(rst),
    .Y(_0967_));
 sky130_fd_sc_hd__inv_2 _3306_ (.A(rst),
    .Y(_0968_));
 sky130_fd_sc_hd__inv_2 _3307_ (.A(rst),
    .Y(_0969_));
 sky130_fd_sc_hd__inv_2 _3308_ (.A(rst),
    .Y(_0970_));
 sky130_fd_sc_hd__inv_2 _3309_ (.A(rst),
    .Y(_0971_));
 sky130_fd_sc_hd__inv_2 _3310_ (.A(rst),
    .Y(_0972_));
 sky130_fd_sc_hd__inv_2 _3311_ (.A(rst),
    .Y(_0973_));
 sky130_fd_sc_hd__inv_2 _3312_ (.A(rst),
    .Y(_0974_));
 sky130_fd_sc_hd__inv_2 _3313_ (.A(rst),
    .Y(_0975_));
 sky130_fd_sc_hd__inv_2 _3314_ (.A(rst),
    .Y(_0976_));
 sky130_fd_sc_hd__inv_2 _3315_ (.A(rst),
    .Y(_0977_));
 sky130_fd_sc_hd__inv_2 _3316_ (.A(rst),
    .Y(_0978_));
 sky130_fd_sc_hd__inv_2 _3317_ (.A(rst),
    .Y(_0979_));
 sky130_fd_sc_hd__inv_2 _3318_ (.A(rst),
    .Y(_0980_));
 sky130_fd_sc_hd__inv_2 _3319_ (.A(rst),
    .Y(_0981_));
 sky130_fd_sc_hd__inv_2 _3320_ (.A(rst),
    .Y(_0982_));
 sky130_fd_sc_hd__inv_2 _3321_ (.A(rst),
    .Y(_0983_));
 sky130_fd_sc_hd__inv_2 _3322_ (.A(rst),
    .Y(_0984_));
 sky130_fd_sc_hd__inv_2 _3323_ (.A(rst),
    .Y(_0985_));
 sky130_fd_sc_hd__inv_2 _3324_ (.A(rst),
    .Y(_0986_));
 sky130_fd_sc_hd__inv_2 _3325_ (.A(rst),
    .Y(_0987_));
 sky130_fd_sc_hd__inv_2 _3326_ (.A(rst),
    .Y(_0988_));
 sky130_fd_sc_hd__inv_2 _3327_ (.A(rst),
    .Y(_0989_));
 sky130_fd_sc_hd__inv_2 _3328_ (.A(rst),
    .Y(_0990_));
 sky130_fd_sc_hd__inv_2 _3329_ (.A(rst),
    .Y(_0991_));
 sky130_fd_sc_hd__inv_2 _3330_ (.A(rst),
    .Y(_0992_));
 sky130_fd_sc_hd__inv_2 _3331_ (.A(rst),
    .Y(_0993_));
 sky130_fd_sc_hd__inv_2 _3332_ (.A(rst),
    .Y(_0994_));
 sky130_fd_sc_hd__inv_2 _3333_ (.A(rst),
    .Y(_0995_));
 sky130_fd_sc_hd__inv_2 _3334_ (.A(rst),
    .Y(_0996_));
 sky130_fd_sc_hd__inv_2 _3335_ (.A(rst),
    .Y(_0997_));
 sky130_fd_sc_hd__inv_2 _3336_ (.A(rst),
    .Y(_0998_));
 sky130_fd_sc_hd__inv_2 _3337_ (.A(rst),
    .Y(_0999_));
 sky130_fd_sc_hd__inv_2 _3338_ (.A(rst),
    .Y(_1000_));
 sky130_fd_sc_hd__inv_2 _3339_ (.A(rst),
    .Y(_1001_));
 sky130_fd_sc_hd__inv_2 _3340_ (.A(rst),
    .Y(_1002_));
 sky130_fd_sc_hd__inv_2 _3341_ (.A(rst),
    .Y(_1003_));
 sky130_fd_sc_hd__inv_2 _3342_ (.A(rst),
    .Y(_1004_));
 sky130_fd_sc_hd__inv_2 _3343_ (.A(rst),
    .Y(_1005_));
 sky130_fd_sc_hd__inv_2 _3344_ (.A(rst),
    .Y(_1006_));
 sky130_fd_sc_hd__inv_2 _3345_ (.A(rst),
    .Y(_1007_));
 sky130_fd_sc_hd__inv_2 _3346_ (.A(rst),
    .Y(_1008_));
 sky130_fd_sc_hd__inv_2 _3347_ (.A(rst),
    .Y(_1009_));
 sky130_fd_sc_hd__inv_2 _3348_ (.A(rst),
    .Y(_1010_));
 sky130_fd_sc_hd__inv_2 _3349_ (.A(rst),
    .Y(_1011_));
 sky130_fd_sc_hd__inv_2 _3350_ (.A(rst),
    .Y(_1012_));
 sky130_fd_sc_hd__inv_2 _3351_ (.A(rst),
    .Y(_1013_));
 sky130_fd_sc_hd__inv_2 _3352_ (.A(rst),
    .Y(_1014_));
 sky130_fd_sc_hd__inv_2 _3353_ (.A(rst),
    .Y(_1015_));
 sky130_fd_sc_hd__inv_2 _3354_ (.A(rst),
    .Y(_1016_));
 sky130_fd_sc_hd__inv_2 _3355_ (.A(rst),
    .Y(_1017_));
 sky130_fd_sc_hd__inv_2 _3356_ (.A(rst),
    .Y(_1018_));
 sky130_fd_sc_hd__inv_2 _3357_ (.A(rst),
    .Y(_1019_));
 sky130_fd_sc_hd__inv_2 _3358_ (.A(rst),
    .Y(_1020_));
 sky130_fd_sc_hd__inv_2 _3359_ (.A(rst),
    .Y(_1021_));
 sky130_fd_sc_hd__inv_2 _3360_ (.A(rst),
    .Y(_1022_));
 sky130_fd_sc_hd__inv_2 _3361_ (.A(rst),
    .Y(_1023_));
 sky130_fd_sc_hd__inv_2 _3362_ (.A(rst),
    .Y(_1024_));
 sky130_fd_sc_hd__inv_2 _3363_ (.A(rst),
    .Y(_1025_));
 sky130_fd_sc_hd__inv_2 _3364_ (.A(rst),
    .Y(_1026_));
 sky130_fd_sc_hd__inv_2 _3365_ (.A(rst),
    .Y(_1027_));
 sky130_fd_sc_hd__inv_2 _3366_ (.A(rst),
    .Y(_1028_));
 sky130_fd_sc_hd__inv_2 _3367_ (.A(rst),
    .Y(_1029_));
 sky130_fd_sc_hd__inv_2 _3368_ (.A(rst),
    .Y(_1030_));
 sky130_fd_sc_hd__inv_2 _3369_ (.A(rst),
    .Y(_1031_));
 sky130_fd_sc_hd__inv_2 _3370_ (.A(rst),
    .Y(_1032_));
 sky130_fd_sc_hd__inv_2 _3371_ (.A(rst),
    .Y(_1033_));
 sky130_fd_sc_hd__inv_2 _3372_ (.A(rst),
    .Y(_1034_));
 sky130_fd_sc_hd__inv_2 _3373_ (.A(rst),
    .Y(_1035_));
 sky130_fd_sc_hd__inv_2 _3374_ (.A(rst),
    .Y(_1036_));
 sky130_fd_sc_hd__inv_2 _3375_ (.A(rst),
    .Y(_1037_));
 sky130_fd_sc_hd__inv_2 _3376_ (.A(rst),
    .Y(_1038_));
 sky130_fd_sc_hd__inv_2 _3377_ (.A(rst),
    .Y(_1039_));
 sky130_fd_sc_hd__inv_2 _3378_ (.A(rst),
    .Y(_1040_));
 sky130_fd_sc_hd__inv_2 _3379_ (.A(rst),
    .Y(_1041_));
 sky130_fd_sc_hd__inv_2 _3380_ (.A(rst),
    .Y(_1042_));
 sky130_fd_sc_hd__inv_2 _3381_ (.A(rst),
    .Y(_1043_));
 sky130_fd_sc_hd__inv_2 _3382_ (.A(rst),
    .Y(_1044_));
 sky130_fd_sc_hd__inv_2 _3383_ (.A(rst),
    .Y(_1045_));
 sky130_fd_sc_hd__inv_2 _3384_ (.A(rst),
    .Y(_1046_));
 sky130_fd_sc_hd__inv_2 _3385_ (.A(rst),
    .Y(_1047_));
 sky130_fd_sc_hd__inv_2 _3386_ (.A(rst),
    .Y(_1048_));
 sky130_fd_sc_hd__inv_2 _3387_ (.A(rst),
    .Y(_1049_));
 sky130_fd_sc_hd__inv_2 _3388_ (.A(rst),
    .Y(_1050_));
 sky130_fd_sc_hd__inv_2 _3389_ (.A(rst),
    .Y(_1051_));
 sky130_fd_sc_hd__inv_2 _3390_ (.A(rst),
    .Y(_1052_));
 sky130_fd_sc_hd__inv_2 _3391_ (.A(rst),
    .Y(_1053_));
 sky130_fd_sc_hd__inv_2 _3392_ (.A(rst),
    .Y(_1054_));
 sky130_fd_sc_hd__inv_2 _3393_ (.A(rst),
    .Y(_1055_));
 sky130_fd_sc_hd__inv_2 _3394_ (.A(rst),
    .Y(_1056_));
 sky130_fd_sc_hd__inv_2 _3395_ (.A(rst),
    .Y(_1057_));
 sky130_fd_sc_hd__inv_2 _3396_ (.A(rst),
    .Y(_1058_));
 sky130_fd_sc_hd__inv_2 _3397_ (.A(rst),
    .Y(_1059_));
 sky130_fd_sc_hd__inv_2 _3398_ (.A(rst),
    .Y(_1060_));
 sky130_fd_sc_hd__inv_2 _3399_ (.A(rst),
    .Y(_1061_));
 sky130_fd_sc_hd__inv_2 _3400_ (.A(rst),
    .Y(_1062_));
 sky130_fd_sc_hd__inv_2 _3401_ (.A(rst),
    .Y(_1063_));
 sky130_fd_sc_hd__inv_2 _3402_ (.A(rst),
    .Y(_1064_));
 sky130_fd_sc_hd__inv_2 _3403_ (.A(rst),
    .Y(_1065_));
 sky130_fd_sc_hd__inv_2 _3404_ (.A(rst),
    .Y(_1066_));
 sky130_fd_sc_hd__inv_2 _3405_ (.A(rst),
    .Y(_1067_));
 sky130_fd_sc_hd__inv_2 _3406_ (.A(rst),
    .Y(_1068_));
 sky130_fd_sc_hd__inv_2 _3407_ (.A(rst),
    .Y(_1069_));
 sky130_fd_sc_hd__inv_2 _3408_ (.A(rst),
    .Y(_1070_));
 sky130_fd_sc_hd__inv_2 _3409_ (.A(rst),
    .Y(_1071_));
 sky130_fd_sc_hd__inv_2 _3410_ (.A(rst),
    .Y(_1072_));
 sky130_fd_sc_hd__inv_2 _3411_ (.A(rst),
    .Y(_1073_));
 sky130_fd_sc_hd__inv_2 _3412_ (.A(rst),
    .Y(_1074_));
 sky130_fd_sc_hd__inv_2 _3413_ (.A(rst),
    .Y(_1075_));
 sky130_fd_sc_hd__inv_2 _3414_ (.A(rst),
    .Y(_1076_));
 sky130_fd_sc_hd__inv_2 _3415_ (.A(rst),
    .Y(_1077_));
 sky130_fd_sc_hd__inv_2 _3416_ (.A(rst),
    .Y(_1078_));
 sky130_fd_sc_hd__inv_2 _3417_ (.A(rst),
    .Y(_1079_));
 sky130_fd_sc_hd__inv_2 _3418_ (.A(rst),
    .Y(_1080_));
 sky130_fd_sc_hd__inv_2 _3419_ (.A(rst),
    .Y(_1081_));
 sky130_fd_sc_hd__inv_2 _3420_ (.A(rst),
    .Y(_1082_));
 sky130_fd_sc_hd__inv_2 _3421_ (.A(rst),
    .Y(_1083_));
 sky130_fd_sc_hd__inv_2 _3422_ (.A(rst),
    .Y(_1084_));
 sky130_fd_sc_hd__inv_2 _3423_ (.A(rst),
    .Y(_1085_));
 sky130_fd_sc_hd__inv_2 _3424_ (.A(rst),
    .Y(_1086_));
 sky130_fd_sc_hd__inv_2 _3425_ (.A(rst),
    .Y(_1087_));
 sky130_fd_sc_hd__inv_2 _3426_ (.A(rst),
    .Y(_1088_));
 sky130_fd_sc_hd__inv_2 _3427_ (.A(rst),
    .Y(_1089_));
 sky130_fd_sc_hd__inv_2 _3428_ (.A(rst),
    .Y(_1090_));
 sky130_fd_sc_hd__inv_2 _3429_ (.A(rst),
    .Y(_1091_));
 sky130_fd_sc_hd__inv_2 _3430_ (.A(rst),
    .Y(_1092_));
 sky130_fd_sc_hd__inv_2 _3431_ (.A(rst),
    .Y(_1093_));
 sky130_fd_sc_hd__inv_2 _3432_ (.A(rst),
    .Y(_1094_));
 sky130_fd_sc_hd__inv_2 _3433_ (.A(rst),
    .Y(_1095_));
 sky130_fd_sc_hd__inv_2 _3434_ (.A(rst),
    .Y(_1096_));
 sky130_fd_sc_hd__inv_2 _3435_ (.A(rst),
    .Y(_1097_));
 sky130_fd_sc_hd__inv_2 _3436_ (.A(rst),
    .Y(_1098_));
 sky130_fd_sc_hd__inv_2 _3437_ (.A(rst),
    .Y(_1099_));
 sky130_fd_sc_hd__inv_2 _3438_ (.A(rst),
    .Y(_1100_));
 sky130_fd_sc_hd__inv_2 _3439_ (.A(rst),
    .Y(_1101_));
 sky130_fd_sc_hd__inv_2 _3440_ (.A(rst),
    .Y(_1102_));
 sky130_fd_sc_hd__inv_2 _3441_ (.A(rst),
    .Y(_1103_));
 sky130_fd_sc_hd__inv_2 _3442_ (.A(rst),
    .Y(_1104_));
 sky130_fd_sc_hd__inv_2 _3443_ (.A(rst),
    .Y(_1105_));
 sky130_fd_sc_hd__inv_2 _3444_ (.A(rst),
    .Y(_1106_));
 sky130_fd_sc_hd__inv_2 _3445_ (.A(rst),
    .Y(_1107_));
 sky130_fd_sc_hd__inv_2 _3446_ (.A(rst),
    .Y(_1108_));
 sky130_fd_sc_hd__inv_2 _3447_ (.A(rst),
    .Y(_1109_));
 sky130_fd_sc_hd__inv_2 _3448_ (.A(rst),
    .Y(_1110_));
 sky130_fd_sc_hd__inv_2 _3449_ (.A(rst),
    .Y(_1111_));
 sky130_fd_sc_hd__inv_2 _3450_ (.A(rst),
    .Y(_1112_));
 sky130_fd_sc_hd__inv_2 _3451_ (.A(rst),
    .Y(_1113_));
 sky130_fd_sc_hd__inv_2 _3452_ (.A(rst),
    .Y(_1114_));
 sky130_fd_sc_hd__inv_2 _3453_ (.A(rst),
    .Y(_1115_));
 sky130_fd_sc_hd__inv_2 _3454_ (.A(rst),
    .Y(_1116_));
 sky130_fd_sc_hd__inv_2 _3455_ (.A(rst),
    .Y(_1117_));
 sky130_fd_sc_hd__inv_2 _3456_ (.A(rst),
    .Y(_1118_));
 sky130_fd_sc_hd__inv_2 _3457_ (.A(rst),
    .Y(_1119_));
 sky130_fd_sc_hd__inv_2 _3458_ (.A(rst),
    .Y(_1120_));
 sky130_fd_sc_hd__inv_2 _3459_ (.A(rst),
    .Y(_1121_));
 sky130_fd_sc_hd__inv_2 _3460_ (.A(rst),
    .Y(_1122_));
 sky130_fd_sc_hd__inv_2 _3461_ (.A(rst),
    .Y(_1123_));
 sky130_fd_sc_hd__inv_2 _3462_ (.A(rst),
    .Y(_1124_));
 sky130_fd_sc_hd__inv_2 _3463_ (.A(rst),
    .Y(_1125_));
 sky130_fd_sc_hd__inv_2 _3464_ (.A(rst),
    .Y(_1126_));
 sky130_fd_sc_hd__inv_2 _3465_ (.A(rst),
    .Y(_1127_));
 sky130_fd_sc_hd__inv_2 _3466_ (.A(rst),
    .Y(_1128_));
 sky130_fd_sc_hd__inv_2 _3467_ (.A(rst),
    .Y(_1129_));
 sky130_fd_sc_hd__inv_2 _3468_ (.A(rst),
    .Y(_1130_));
 sky130_fd_sc_hd__inv_2 _3469_ (.A(rst),
    .Y(_1131_));
 sky130_fd_sc_hd__inv_2 _3470_ (.A(rst),
    .Y(_1132_));
 sky130_fd_sc_hd__inv_2 _3471_ (.A(rst),
    .Y(_1133_));
 sky130_fd_sc_hd__inv_2 _3472_ (.A(rst),
    .Y(_1134_));
 sky130_fd_sc_hd__inv_2 _3473_ (.A(rst),
    .Y(_1135_));
 sky130_fd_sc_hd__inv_2 _3474_ (.A(rst),
    .Y(_1136_));
 sky130_fd_sc_hd__inv_2 _3475_ (.A(rst),
    .Y(_1137_));
 sky130_fd_sc_hd__inv_2 _3476_ (.A(rst),
    .Y(_1138_));
 sky130_fd_sc_hd__inv_2 _3477_ (.A(rst),
    .Y(_1139_));
 sky130_fd_sc_hd__inv_2 _3478_ (.A(rst),
    .Y(_1140_));
 sky130_fd_sc_hd__inv_2 _3479_ (.A(rst),
    .Y(_1141_));
 sky130_fd_sc_hd__inv_2 _3480_ (.A(rst),
    .Y(_1142_));
 sky130_fd_sc_hd__inv_2 _3481_ (.A(rst),
    .Y(_1143_));
 sky130_fd_sc_hd__inv_2 _3482_ (.A(rst),
    .Y(_1144_));
 sky130_fd_sc_hd__inv_2 _3483_ (.A(rst),
    .Y(_1145_));
 sky130_fd_sc_hd__inv_2 _3484_ (.A(rst),
    .Y(_1146_));
 sky130_fd_sc_hd__inv_2 _3485_ (.A(rst),
    .Y(_1147_));
 sky130_fd_sc_hd__inv_2 _3486_ (.A(rst),
    .Y(_1148_));
 sky130_fd_sc_hd__inv_2 _3487_ (.A(rst),
    .Y(_1149_));
 sky130_fd_sc_hd__inv_2 _3488_ (.A(rst),
    .Y(_1150_));
 sky130_fd_sc_hd__inv_2 _3489_ (.A(rst),
    .Y(_1151_));
 sky130_fd_sc_hd__inv_2 _3490_ (.A(rst),
    .Y(_1152_));
 sky130_fd_sc_hd__inv_2 _3491_ (.A(rst),
    .Y(_1153_));
 sky130_fd_sc_hd__inv_2 _3492_ (.A(rst),
    .Y(_1154_));
 sky130_fd_sc_hd__inv_2 _3493_ (.A(rst),
    .Y(_1155_));
 sky130_fd_sc_hd__inv_2 _3494_ (.A(rst),
    .Y(_1156_));
 sky130_fd_sc_hd__inv_2 _3495_ (.A(rst),
    .Y(_1157_));
 sky130_fd_sc_hd__inv_2 _3496_ (.A(rst),
    .Y(_1158_));
 sky130_fd_sc_hd__inv_2 _3497_ (.A(rst),
    .Y(_1159_));
 sky130_fd_sc_hd__inv_2 _3498_ (.A(rst),
    .Y(_1160_));
 sky130_fd_sc_hd__inv_2 _3499_ (.A(rst),
    .Y(_1161_));
 sky130_fd_sc_hd__inv_2 _3500_ (.A(rst),
    .Y(_1162_));
 sky130_fd_sc_hd__inv_2 _3501_ (.A(rst),
    .Y(_1163_));
 sky130_fd_sc_hd__inv_2 _3502_ (.A(rst),
    .Y(_1164_));
 sky130_fd_sc_hd__inv_2 _3503_ (.A(rst),
    .Y(_1165_));
 sky130_fd_sc_hd__inv_2 _3504_ (.A(rst),
    .Y(_1166_));
 sky130_fd_sc_hd__inv_2 _3505_ (.A(rst),
    .Y(_1167_));
 sky130_fd_sc_hd__inv_2 _3506_ (.A(rst),
    .Y(_1168_));
 sky130_fd_sc_hd__inv_2 _3507_ (.A(rst),
    .Y(_1169_));
 sky130_fd_sc_hd__inv_2 _3508_ (.A(rst),
    .Y(_1170_));
 sky130_fd_sc_hd__inv_2 _3509_ (.A(rst),
    .Y(_1171_));
 sky130_fd_sc_hd__inv_2 _3510_ (.A(rst),
    .Y(_1172_));
 sky130_fd_sc_hd__inv_2 _3511_ (.A(rst),
    .Y(_1173_));
 sky130_fd_sc_hd__inv_2 _3512_ (.A(rst),
    .Y(_1174_));
 sky130_fd_sc_hd__inv_2 _3513_ (.A(rst),
    .Y(_1175_));
 sky130_fd_sc_hd__inv_2 _3514_ (.A(rst),
    .Y(_1176_));
 sky130_fd_sc_hd__inv_2 _3515_ (.A(rst),
    .Y(_1177_));
 sky130_fd_sc_hd__inv_2 _3516_ (.A(rst),
    .Y(_1178_));
 sky130_fd_sc_hd__inv_2 _3517_ (.A(rst),
    .Y(_1179_));
 sky130_fd_sc_hd__inv_2 _3518_ (.A(rst),
    .Y(_1180_));
 sky130_fd_sc_hd__inv_2 _3519_ (.A(rst),
    .Y(_1181_));
 sky130_fd_sc_hd__inv_2 _3520_ (.A(rst),
    .Y(_1182_));
 sky130_fd_sc_hd__inv_2 _3521_ (.A(rst),
    .Y(_1183_));
 sky130_fd_sc_hd__inv_2 _3522_ (.A(rst),
    .Y(_1184_));
 sky130_fd_sc_hd__inv_2 _3523_ (.A(rst),
    .Y(_1185_));
 sky130_fd_sc_hd__inv_2 _3524_ (.A(rst),
    .Y(_1186_));
 sky130_fd_sc_hd__inv_2 _3525_ (.A(rst),
    .Y(_1187_));
 sky130_fd_sc_hd__inv_2 _3526_ (.A(rst),
    .Y(_1188_));
 sky130_fd_sc_hd__inv_2 _3527_ (.A(rst),
    .Y(_1189_));
 sky130_fd_sc_hd__inv_2 _3528_ (.A(rst),
    .Y(_1190_));
 sky130_fd_sc_hd__inv_2 _3529_ (.A(rst),
    .Y(_1191_));
 sky130_fd_sc_hd__inv_2 _3530_ (.A(rst),
    .Y(_1192_));
 sky130_fd_sc_hd__inv_2 _3531_ (.A(rst),
    .Y(_1193_));
 sky130_fd_sc_hd__inv_2 _3532_ (.A(rst),
    .Y(_1194_));
 sky130_fd_sc_hd__inv_2 _3533_ (.A(rst),
    .Y(_1195_));
 sky130_fd_sc_hd__inv_2 _3534_ (.A(rst),
    .Y(_1196_));
 sky130_fd_sc_hd__inv_2 _3535_ (.A(rst),
    .Y(_1197_));
 sky130_fd_sc_hd__inv_2 _3536_ (.A(rst),
    .Y(_1198_));
 sky130_fd_sc_hd__inv_2 _3537_ (.A(rst),
    .Y(_1199_));
 sky130_fd_sc_hd__inv_2 _3538_ (.A(rst),
    .Y(_1200_));
 sky130_fd_sc_hd__inv_2 _3539_ (.A(rst),
    .Y(_1201_));
 sky130_fd_sc_hd__inv_2 _3540_ (.A(rst),
    .Y(_1202_));
 sky130_fd_sc_hd__inv_2 _3541_ (.A(rst),
    .Y(_1203_));
 sky130_fd_sc_hd__inv_2 _3542_ (.A(rst),
    .Y(_1204_));
 sky130_fd_sc_hd__inv_2 _3543_ (.A(rst),
    .Y(_1205_));
 sky130_fd_sc_hd__inv_2 _3544_ (.A(rst),
    .Y(_1206_));
 sky130_fd_sc_hd__inv_2 _3545_ (.A(rst),
    .Y(_1207_));
 sky130_fd_sc_hd__inv_2 _3546_ (.A(rst),
    .Y(_1208_));
 sky130_fd_sc_hd__inv_2 _3547_ (.A(rst),
    .Y(_1209_));
 sky130_fd_sc_hd__inv_2 _3548_ (.A(rst),
    .Y(_1210_));
 sky130_fd_sc_hd__inv_2 _3549_ (.A(rst),
    .Y(_1211_));
 sky130_fd_sc_hd__inv_2 _3550_ (.A(rst),
    .Y(_1212_));
 sky130_fd_sc_hd__inv_2 _3551_ (.A(rst),
    .Y(_1213_));
 sky130_fd_sc_hd__inv_2 _3552_ (.A(rst),
    .Y(_1214_));
 sky130_fd_sc_hd__inv_2 _3553_ (.A(rst),
    .Y(_1215_));
 sky130_fd_sc_hd__inv_2 _3554_ (.A(rst),
    .Y(_1216_));
 sky130_fd_sc_hd__inv_2 _3555_ (.A(rst),
    .Y(_1217_));
 sky130_fd_sc_hd__inv_2 _3556_ (.A(rst),
    .Y(_1218_));
 sky130_fd_sc_hd__inv_2 _3557_ (.A(rst),
    .Y(_1219_));
 sky130_fd_sc_hd__inv_2 _3558_ (.A(rst),
    .Y(_1220_));
 sky130_fd_sc_hd__inv_2 _3559_ (.A(rst),
    .Y(_1221_));
 sky130_fd_sc_hd__inv_2 _3560_ (.A(rst),
    .Y(_1222_));
 sky130_fd_sc_hd__inv_2 _3561_ (.A(rst),
    .Y(_1223_));
 sky130_fd_sc_hd__inv_2 _3562_ (.A(rst),
    .Y(_1224_));
 sky130_fd_sc_hd__inv_2 _3563_ (.A(rst),
    .Y(_1225_));
 sky130_fd_sc_hd__inv_2 _3564_ (.A(rst),
    .Y(_1226_));
 sky130_fd_sc_hd__inv_2 _3565_ (.A(rst),
    .Y(_1227_));
 sky130_fd_sc_hd__inv_2 _3566_ (.A(rst),
    .Y(_1228_));
 sky130_fd_sc_hd__inv_2 _3567_ (.A(rst),
    .Y(_1229_));
 sky130_fd_sc_hd__inv_2 _3568_ (.A(rst),
    .Y(_1230_));
 sky130_fd_sc_hd__inv_2 _3569_ (.A(rst),
    .Y(_1231_));
 sky130_fd_sc_hd__inv_2 _3570_ (.A(rst),
    .Y(_1232_));
 sky130_fd_sc_hd__inv_2 _3571_ (.A(rst),
    .Y(_1233_));
 sky130_fd_sc_hd__inv_2 _3572_ (.A(rst),
    .Y(_1234_));
 sky130_fd_sc_hd__inv_2 _3573_ (.A(rst),
    .Y(_1235_));
 sky130_fd_sc_hd__inv_2 _3574_ (.A(rst),
    .Y(_1236_));
 sky130_fd_sc_hd__inv_2 _3575_ (.A(rst),
    .Y(_1237_));
 sky130_fd_sc_hd__inv_2 _3576_ (.A(rst),
    .Y(_1238_));
 sky130_fd_sc_hd__inv_2 _3577_ (.A(rst),
    .Y(_1239_));
 sky130_fd_sc_hd__inv_2 _3578_ (.A(rst),
    .Y(_1240_));
 sky130_fd_sc_hd__inv_2 _3579_ (.A(rst),
    .Y(_1241_));
 sky130_fd_sc_hd__inv_2 _3580_ (.A(rst),
    .Y(_1242_));
 sky130_fd_sc_hd__inv_2 _3581_ (.A(rst),
    .Y(_1243_));
 sky130_fd_sc_hd__inv_2 _3582_ (.A(rst),
    .Y(_1244_));
 sky130_fd_sc_hd__inv_2 _3583_ (.A(rst),
    .Y(_1245_));
 sky130_fd_sc_hd__inv_2 _3584_ (.A(rst),
    .Y(_1246_));
 sky130_fd_sc_hd__inv_2 _3585_ (.A(rst),
    .Y(_1247_));
 sky130_fd_sc_hd__inv_2 _3586_ (.A(rst),
    .Y(_1248_));
 sky130_fd_sc_hd__inv_2 _3587_ (.A(rst),
    .Y(_1249_));
 sky130_fd_sc_hd__inv_2 _3588_ (.A(rst),
    .Y(_1250_));
 sky130_fd_sc_hd__inv_2 _3589_ (.A(rst),
    .Y(_1251_));
 sky130_fd_sc_hd__inv_2 _3590_ (.A(rst),
    .Y(_1252_));
 sky130_fd_sc_hd__inv_2 _3591_ (.A(rst),
    .Y(_1253_));
 sky130_fd_sc_hd__inv_2 _3592_ (.A(rst),
    .Y(_1254_));
 sky130_fd_sc_hd__inv_2 _3593_ (.A(rst),
    .Y(_1255_));
 sky130_fd_sc_hd__inv_2 _3594_ (.A(rst),
    .Y(_1256_));
 sky130_fd_sc_hd__inv_2 _3595_ (.A(rst),
    .Y(_1257_));
 sky130_fd_sc_hd__inv_2 _3596_ (.A(rst),
    .Y(_1258_));
 sky130_fd_sc_hd__inv_2 _3597_ (.A(rst),
    .Y(_1259_));
 sky130_fd_sc_hd__inv_2 _3598_ (.A(rst),
    .Y(_1260_));
 sky130_fd_sc_hd__inv_2 _3599_ (.A(rst),
    .Y(_1261_));
 sky130_fd_sc_hd__inv_2 _3600_ (.A(rst),
    .Y(_1262_));
 sky130_fd_sc_hd__inv_2 _3601_ (.A(rst),
    .Y(_1263_));
 sky130_fd_sc_hd__inv_2 _3602_ (.A(rst),
    .Y(_1264_));
 sky130_fd_sc_hd__inv_2 _3603_ (.A(rst),
    .Y(_1265_));
 sky130_fd_sc_hd__inv_2 _3604_ (.A(rst),
    .Y(_1266_));
 sky130_fd_sc_hd__inv_2 _3605_ (.A(rst),
    .Y(_1267_));
 sky130_fd_sc_hd__inv_2 _3606_ (.A(rst),
    .Y(_1268_));
 sky130_fd_sc_hd__inv_2 _3607_ (.A(rst),
    .Y(_1269_));
 sky130_fd_sc_hd__inv_2 _3608_ (.A(rst),
    .Y(_1270_));
 sky130_fd_sc_hd__inv_2 _3609_ (.A(rst),
    .Y(_1271_));
 sky130_fd_sc_hd__inv_2 _3610_ (.A(rst),
    .Y(_1272_));
 sky130_fd_sc_hd__inv_2 _3611_ (.A(rst),
    .Y(_1273_));
 sky130_fd_sc_hd__inv_2 _3612_ (.A(rst),
    .Y(_1274_));
 sky130_fd_sc_hd__inv_2 _3613_ (.A(rst),
    .Y(_1275_));
 sky130_fd_sc_hd__inv_2 _3614_ (.A(rst),
    .Y(_1276_));
 sky130_fd_sc_hd__inv_2 _3615_ (.A(rst),
    .Y(_1277_));
 sky130_fd_sc_hd__inv_2 _3616_ (.A(rst),
    .Y(_1278_));
 sky130_fd_sc_hd__inv_2 _3617_ (.A(rst),
    .Y(_1279_));
 sky130_fd_sc_hd__inv_2 _3618_ (.A(rst),
    .Y(_1280_));
 sky130_fd_sc_hd__inv_2 _3619_ (.A(rst),
    .Y(_1281_));
 sky130_fd_sc_hd__inv_2 _3620_ (.A(rst),
    .Y(_1282_));
 sky130_fd_sc_hd__inv_2 _3621_ (.A(rst),
    .Y(_1283_));
 sky130_fd_sc_hd__inv_2 _3622_ (.A(rst),
    .Y(_1284_));
 sky130_fd_sc_hd__inv_2 _3623_ (.A(rst),
    .Y(_1285_));
 sky130_fd_sc_hd__inv_2 _3624_ (.A(rst),
    .Y(_1286_));
 sky130_fd_sc_hd__inv_2 _3625_ (.A(rst),
    .Y(_1287_));
 sky130_fd_sc_hd__inv_2 _3626_ (.A(rst),
    .Y(_1288_));
 sky130_fd_sc_hd__inv_2 _3627_ (.A(rst),
    .Y(_1289_));
 sky130_fd_sc_hd__inv_2 _3628_ (.A(rst),
    .Y(_1290_));
 sky130_fd_sc_hd__inv_2 _3629_ (.A(rst),
    .Y(_1291_));
 sky130_fd_sc_hd__inv_2 _3630_ (.A(rst),
    .Y(_1292_));
 sky130_fd_sc_hd__inv_2 _3631_ (.A(rst),
    .Y(_1293_));
 sky130_fd_sc_hd__inv_2 _3632_ (.A(rst),
    .Y(_1294_));
 sky130_fd_sc_hd__inv_2 _3633_ (.A(rst),
    .Y(_1295_));
 sky130_fd_sc_hd__inv_2 _3634_ (.A(rst),
    .Y(_1296_));
 sky130_fd_sc_hd__inv_2 _3635_ (.A(rst),
    .Y(_1297_));
 sky130_fd_sc_hd__inv_2 _3636_ (.A(rst),
    .Y(_1298_));
 sky130_fd_sc_hd__inv_2 _3637_ (.A(rst),
    .Y(_1299_));
 sky130_fd_sc_hd__inv_2 _3638_ (.A(rst),
    .Y(_1300_));
 sky130_fd_sc_hd__inv_2 _3639_ (.A(rst),
    .Y(_1301_));
 sky130_fd_sc_hd__inv_2 _3640_ (.A(rst),
    .Y(_1302_));
 sky130_fd_sc_hd__inv_2 _3641_ (.A(rst),
    .Y(_1303_));
 sky130_fd_sc_hd__inv_2 _3642_ (.A(rst),
    .Y(_1304_));
 sky130_fd_sc_hd__inv_2 _3643_ (.A(rst),
    .Y(_1305_));
 sky130_fd_sc_hd__inv_2 _3644_ (.A(rst),
    .Y(_1306_));
 sky130_fd_sc_hd__inv_2 _3645_ (.A(rst),
    .Y(_1307_));
 sky130_fd_sc_hd__inv_2 _3646_ (.A(rst),
    .Y(_1308_));
 sky130_fd_sc_hd__inv_2 _3647_ (.A(rst),
    .Y(_1309_));
 sky130_fd_sc_hd__inv_2 _3648_ (.A(rst),
    .Y(_1310_));
 sky130_fd_sc_hd__inv_2 _3649_ (.A(rst),
    .Y(_1311_));
 sky130_fd_sc_hd__inv_2 _3650_ (.A(rst),
    .Y(_1312_));
 sky130_fd_sc_hd__inv_2 _3651_ (.A(rst),
    .Y(_1313_));
 sky130_fd_sc_hd__inv_2 _3652_ (.A(rst),
    .Y(_1314_));
 sky130_fd_sc_hd__inv_2 _3653_ (.A(rst),
    .Y(_1315_));
 sky130_fd_sc_hd__inv_2 _3654_ (.A(rst),
    .Y(_1316_));
 sky130_fd_sc_hd__inv_2 _3655_ (.A(rst),
    .Y(_1317_));
 sky130_fd_sc_hd__inv_2 _3656_ (.A(rst),
    .Y(_1318_));
 sky130_fd_sc_hd__inv_2 _3657_ (.A(rst),
    .Y(_1319_));
 sky130_fd_sc_hd__inv_2 _3658_ (.A(rst),
    .Y(_1320_));
 sky130_fd_sc_hd__inv_2 _3659_ (.A(rst),
    .Y(_1321_));
 sky130_fd_sc_hd__inv_2 _3660_ (.A(rst),
    .Y(_1322_));
 sky130_fd_sc_hd__inv_2 _3661_ (.A(rst),
    .Y(_1323_));
 sky130_fd_sc_hd__inv_2 _3662_ (.A(rst),
    .Y(_1324_));
 sky130_fd_sc_hd__inv_2 _3663_ (.A(rst),
    .Y(_1325_));
 sky130_fd_sc_hd__inv_2 _3664_ (.A(rst),
    .Y(_1326_));
 sky130_fd_sc_hd__inv_2 _3665_ (.A(rst),
    .Y(_1327_));
 sky130_fd_sc_hd__inv_2 _3666_ (.A(rst),
    .Y(_1328_));
 sky130_fd_sc_hd__inv_2 _3667_ (.A(rst),
    .Y(_1329_));
 sky130_fd_sc_hd__inv_2 _3668_ (.A(rst),
    .Y(_1330_));
 sky130_fd_sc_hd__inv_2 _3669_ (.A(rst),
    .Y(_1331_));
 sky130_fd_sc_hd__inv_2 _3670_ (.A(rst),
    .Y(_1332_));
 sky130_fd_sc_hd__inv_2 _3671_ (.A(rst),
    .Y(_1333_));
 sky130_fd_sc_hd__inv_2 _3672_ (.A(rst),
    .Y(_1334_));
 sky130_fd_sc_hd__inv_2 _3673_ (.A(rst),
    .Y(_1335_));
 sky130_fd_sc_hd__inv_2 _3674_ (.A(rst),
    .Y(_1336_));
 sky130_fd_sc_hd__inv_2 _3675_ (.A(rst),
    .Y(_1337_));
 sky130_fd_sc_hd__inv_2 _3676_ (.A(rst),
    .Y(_1338_));
 sky130_fd_sc_hd__inv_2 _3677_ (.A(rst),
    .Y(_1339_));
 sky130_fd_sc_hd__inv_2 _3678_ (.A(rst),
    .Y(_1340_));
 sky130_fd_sc_hd__inv_2 _3679_ (.A(rst),
    .Y(_1341_));
 sky130_fd_sc_hd__inv_2 _3680_ (.A(rst),
    .Y(_1342_));
 sky130_fd_sc_hd__inv_2 _3681_ (.A(rst),
    .Y(_1343_));
 sky130_fd_sc_hd__inv_2 _3682_ (.A(rst),
    .Y(_1344_));
 sky130_fd_sc_hd__inv_2 _3683_ (.A(rst),
    .Y(_1345_));
 sky130_fd_sc_hd__inv_2 _3684_ (.A(out_data_flat[26]),
    .Y(_1410_));
 sky130_fd_sc_hd__inv_2 _3685_ (.A(out_data_flat[24]),
    .Y(_1411_));
 sky130_fd_sc_hd__inv_2 _3686_ (.A(out_data_flat[14]),
    .Y(_1412_));
 sky130_fd_sc_hd__inv_2 _3687_ (.A(out_data_flat[9]),
    .Y(_1413_));
 sky130_fd_sc_hd__inv_2 _3688_ (.A(out_data_flat[8]),
    .Y(_1414_));
 sky130_fd_sc_hd__inv_2 _3689_ (.A(out_data_flat[4]),
    .Y(_1415_));
 sky130_fd_sc_hd__inv_2 _3690_ (.A(out_data_flat[1]),
    .Y(_1416_));
 sky130_fd_sc_hd__inv_2 _3691_ (.A(out_data_flat[0]),
    .Y(_1417_));
 sky130_fd_sc_hd__inv_2 _3692_ (.A(out_data_flat[254]),
    .Y(_1418_));
 sky130_fd_sc_hd__inv_2 _3693_ (.A(out_data_flat[251]),
    .Y(_1419_));
 sky130_fd_sc_hd__inv_2 _3694_ (.A(out_data_flat[250]),
    .Y(_1420_));
 sky130_fd_sc_hd__inv_2 _3695_ (.A(out_data_flat[249]),
    .Y(_1421_));
 sky130_fd_sc_hd__inv_2 _3696_ (.A(out_data_flat[244]),
    .Y(_1422_));
 sky130_fd_sc_hd__inv_2 _3697_ (.A(out_data_flat[241]),
    .Y(_1423_));
 sky130_fd_sc_hd__inv_2 _3698_ (.A(out_data_flat[239]),
    .Y(_1424_));
 sky130_fd_sc_hd__inv_2 _3699_ (.A(out_data_flat[238]),
    .Y(_1425_));
 sky130_fd_sc_hd__inv_2 _3700_ (.A(out_data_flat[237]),
    .Y(_1426_));
 sky130_fd_sc_hd__inv_2 _3701_ (.A(out_data_flat[236]),
    .Y(_1427_));
 sky130_fd_sc_hd__inv_2 _3702_ (.A(\gen_pe[1].pe_inst.sel ),
    .Y(_1428_));
 sky130_fd_sc_hd__inv_2 _3703_ (.A(out_data_flat[63]),
    .Y(_1429_));
 sky130_fd_sc_hd__inv_2 _3704_ (.A(out_data_flat[62]),
    .Y(_1430_));
 sky130_fd_sc_hd__inv_2 _3705_ (.A(out_data_flat[61]),
    .Y(_1431_));
 sky130_fd_sc_hd__inv_2 _3706_ (.A(out_data_flat[60]),
    .Y(_1432_));
 sky130_fd_sc_hd__inv_2 _3707_ (.A(out_data_flat[57]),
    .Y(_1433_));
 sky130_fd_sc_hd__inv_2 _3708_ (.A(out_data_flat[55]),
    .Y(_1434_));
 sky130_fd_sc_hd__inv_2 _3709_ (.A(out_data_flat[54]),
    .Y(_1435_));
 sky130_fd_sc_hd__inv_2 _3710_ (.A(out_data_flat[53]),
    .Y(_1436_));
 sky130_fd_sc_hd__inv_2 _3711_ (.A(out_data_flat[52]),
    .Y(_1437_));
 sky130_fd_sc_hd__inv_2 _3712_ (.A(out_data_flat[51]),
    .Y(_1438_));
 sky130_fd_sc_hd__inv_2 _3713_ (.A(out_data_flat[50]),
    .Y(_1439_));
 sky130_fd_sc_hd__inv_2 _3714_ (.A(out_data_flat[49]),
    .Y(_1440_));
 sky130_fd_sc_hd__inv_2 _3715_ (.A(out_data_flat[48]),
    .Y(_1441_));
 sky130_fd_sc_hd__inv_2 _3716_ (.A(out_data_flat[47]),
    .Y(_1442_));
 sky130_fd_sc_hd__inv_2 _3717_ (.A(out_data_flat[45]),
    .Y(_1443_));
 sky130_fd_sc_hd__inv_2 _3718_ (.A(out_data_flat[44]),
    .Y(_1444_));
 sky130_fd_sc_hd__inv_2 _3719_ (.A(out_data_flat[43]),
    .Y(_1445_));
 sky130_fd_sc_hd__inv_2 _3720_ (.A(out_data_flat[42]),
    .Y(_1446_));
 sky130_fd_sc_hd__inv_2 _3721_ (.A(out_data_flat[37]),
    .Y(_1447_));
 sky130_fd_sc_hd__inv_2 _3722_ (.A(out_data_flat[34]),
    .Y(_1448_));
 sky130_fd_sc_hd__inv_2 _3723_ (.A(out_data_flat[223]),
    .Y(_1449_));
 sky130_fd_sc_hd__inv_2 _3724_ (.A(out_data_flat[222]),
    .Y(_1450_));
 sky130_fd_sc_hd__inv_2 _3725_ (.A(out_data_flat[221]),
    .Y(_1451_));
 sky130_fd_sc_hd__inv_2 _3726_ (.A(out_data_flat[220]),
    .Y(_1452_));
 sky130_fd_sc_hd__inv_2 _3727_ (.A(out_data_flat[216]),
    .Y(_1453_));
 sky130_fd_sc_hd__inv_2 _3728_ (.A(out_data_flat[213]),
    .Y(_1454_));
 sky130_fd_sc_hd__inv_2 _3729_ (.A(out_data_flat[211]),
    .Y(_1455_));
 sky130_fd_sc_hd__inv_2 _3730_ (.A(out_data_flat[210]),
    .Y(_1456_));
 sky130_fd_sc_hd__inv_2 _3731_ (.A(out_data_flat[208]),
    .Y(_1457_));
 sky130_fd_sc_hd__inv_2 _3732_ (.A(out_data_flat[204]),
    .Y(_1458_));
 sky130_fd_sc_hd__inv_2 _3733_ (.A(out_data_flat[203]),
    .Y(_1459_));
 sky130_fd_sc_hd__inv_2 _3734_ (.A(out_data_flat[202]),
    .Y(_1460_));
 sky130_fd_sc_hd__inv_2 _3735_ (.A(out_data_flat[197]),
    .Y(_1461_));
 sky130_fd_sc_hd__inv_2 _3736_ (.A(out_data_flat[196]),
    .Y(_1462_));
 sky130_fd_sc_hd__inv_2 _3737_ (.A(out_data_flat[195]),
    .Y(_1463_));
 sky130_fd_sc_hd__inv_2 _3738_ (.A(out_data_flat[194]),
    .Y(_1464_));
 sky130_fd_sc_hd__inv_2 _3739_ (.A(out_data_flat[95]),
    .Y(_1465_));
 sky130_fd_sc_hd__inv_2 _3740_ (.A(out_data_flat[94]),
    .Y(_1466_));
 sky130_fd_sc_hd__inv_2 _3741_ (.A(out_data_flat[93]),
    .Y(_1467_));
 sky130_fd_sc_hd__inv_2 _3742_ (.A(out_data_flat[92]),
    .Y(_1468_));
 sky130_fd_sc_hd__inv_2 _3743_ (.A(out_data_flat[91]),
    .Y(_1469_));
 sky130_fd_sc_hd__inv_2 _3744_ (.A(out_data_flat[90]),
    .Y(_1470_));
 sky130_fd_sc_hd__inv_2 _3745_ (.A(out_data_flat[89]),
    .Y(_1471_));
 sky130_fd_sc_hd__inv_2 _3746_ (.A(out_data_flat[88]),
    .Y(_1472_));
 sky130_fd_sc_hd__inv_2 _3747_ (.A(out_data_flat[81]),
    .Y(_1473_));
 sky130_fd_sc_hd__inv_2 _3748_ (.A(out_data_flat[80]),
    .Y(_1474_));
 sky130_fd_sc_hd__inv_2 _3749_ (.A(out_data_flat[78]),
    .Y(_1475_));
 sky130_fd_sc_hd__inv_2 _3750_ (.A(out_data_flat[73]),
    .Y(_1476_));
 sky130_fd_sc_hd__inv_2 _3751_ (.A(out_data_flat[72]),
    .Y(_1477_));
 sky130_fd_sc_hd__inv_2 _3752_ (.A(out_data_flat[71]),
    .Y(_1478_));
 sky130_fd_sc_hd__inv_2 _3753_ (.A(out_data_flat[70]),
    .Y(_1479_));
 sky130_fd_sc_hd__inv_2 _3754_ (.A(out_data_flat[69]),
    .Y(_1480_));
 sky130_fd_sc_hd__inv_2 _3755_ (.A(out_data_flat[68]),
    .Y(_1481_));
 sky130_fd_sc_hd__inv_2 _3756_ (.A(out_data_flat[67]),
    .Y(_1482_));
 sky130_fd_sc_hd__inv_2 _3757_ (.A(out_data_flat[66]),
    .Y(_1483_));
 sky130_fd_sc_hd__inv_2 _3758_ (.A(out_data_flat[65]),
    .Y(_1484_));
 sky130_fd_sc_hd__inv_2 _3759_ (.A(out_data_flat[64]),
    .Y(_1485_));
 sky130_fd_sc_hd__inv_2 _3760_ (.A(out_data_flat[127]),
    .Y(_1486_));
 sky130_fd_sc_hd__inv_2 _3761_ (.A(out_data_flat[126]),
    .Y(_1487_));
 sky130_fd_sc_hd__inv_2 _3762_ (.A(out_data_flat[125]),
    .Y(_1488_));
 sky130_fd_sc_hd__inv_2 _3763_ (.A(out_data_flat[124]),
    .Y(_1489_));
 sky130_fd_sc_hd__inv_2 _3764_ (.A(out_data_flat[123]),
    .Y(_1490_));
 sky130_fd_sc_hd__inv_2 _3765_ (.A(out_data_flat[122]),
    .Y(_1491_));
 sky130_fd_sc_hd__inv_2 _3766_ (.A(out_data_flat[121]),
    .Y(_1492_));
 sky130_fd_sc_hd__inv_2 _3767_ (.A(out_data_flat[120]),
    .Y(_1493_));
 sky130_fd_sc_hd__inv_2 _3768_ (.A(out_data_flat[119]),
    .Y(_1494_));
 sky130_fd_sc_hd__inv_2 _3769_ (.A(out_data_flat[118]),
    .Y(_1495_));
 sky130_fd_sc_hd__inv_2 _3770_ (.A(out_data_flat[117]),
    .Y(_1496_));
 sky130_fd_sc_hd__inv_2 _3771_ (.A(out_data_flat[116]),
    .Y(_1497_));
 sky130_fd_sc_hd__inv_2 _3772_ (.A(out_data_flat[115]),
    .Y(_1498_));
 sky130_fd_sc_hd__inv_2 _3773_ (.A(out_data_flat[114]),
    .Y(_1499_));
 sky130_fd_sc_hd__inv_2 _3774_ (.A(out_data_flat[113]),
    .Y(_1500_));
 sky130_fd_sc_hd__inv_2 _3775_ (.A(out_data_flat[112]),
    .Y(_1501_));
 sky130_fd_sc_hd__inv_2 _3776_ (.A(out_data_flat[111]),
    .Y(_1502_));
 sky130_fd_sc_hd__inv_2 _3777_ (.A(out_data_flat[101]),
    .Y(_1503_));
 sky130_fd_sc_hd__inv_2 _3778_ (.A(out_data_flat[190]),
    .Y(_1504_));
 sky130_fd_sc_hd__inv_2 _3779_ (.A(out_data_flat[189]),
    .Y(_1505_));
 sky130_fd_sc_hd__inv_2 _3780_ (.A(out_data_flat[188]),
    .Y(_1506_));
 sky130_fd_sc_hd__inv_2 _3781_ (.A(out_data_flat[185]),
    .Y(_1507_));
 sky130_fd_sc_hd__inv_2 _3782_ (.A(out_data_flat[184]),
    .Y(_1508_));
 sky130_fd_sc_hd__inv_2 _3783_ (.A(out_data_flat[183]),
    .Y(_1509_));
 sky130_fd_sc_hd__inv_2 _3784_ (.A(out_data_flat[182]),
    .Y(_1510_));
 sky130_fd_sc_hd__inv_2 _3785_ (.A(out_data_flat[181]),
    .Y(_1511_));
 sky130_fd_sc_hd__inv_2 _3786_ (.A(out_data_flat[180]),
    .Y(_1512_));
 sky130_fd_sc_hd__inv_2 _3787_ (.A(out_data_flat[177]),
    .Y(_1513_));
 sky130_fd_sc_hd__inv_2 _3788_ (.A(out_data_flat[176]),
    .Y(_1514_));
 sky130_fd_sc_hd__inv_2 _3789_ (.A(out_data_flat[173]),
    .Y(_1515_));
 sky130_fd_sc_hd__inv_2 _3790_ (.A(out_data_flat[169]),
    .Y(_1516_));
 sky130_fd_sc_hd__inv_2 _3791_ (.A(out_data_flat[168]),
    .Y(_1517_));
 sky130_fd_sc_hd__inv_2 _3792_ (.A(out_data_flat[165]),
    .Y(_1518_));
 sky130_fd_sc_hd__inv_2 _3793_ (.A(out_data_flat[162]),
    .Y(_1519_));
 sky130_fd_sc_hd__inv_2 _3794_ (.A(out_data_flat[160]),
    .Y(_1520_));
 sky130_fd_sc_hd__inv_2 _3795_ (.A(out_data_flat[159]),
    .Y(_1521_));
 sky130_fd_sc_hd__inv_2 _3796_ (.A(out_data_flat[156]),
    .Y(_1522_));
 sky130_fd_sc_hd__inv_2 _3797_ (.A(out_data_flat[155]),
    .Y(_1523_));
 sky130_fd_sc_hd__inv_2 _3798_ (.A(out_data_flat[152]),
    .Y(_1524_));
 sky130_fd_sc_hd__inv_2 _3799_ (.A(out_data_flat[151]),
    .Y(_1525_));
 sky130_fd_sc_hd__inv_2 _3800_ (.A(out_data_flat[148]),
    .Y(_1526_));
 sky130_fd_sc_hd__inv_2 _3801_ (.A(out_data_flat[145]),
    .Y(_1527_));
 sky130_fd_sc_hd__inv_2 _3802_ (.A(out_data_flat[144]),
    .Y(_1528_));
 sky130_fd_sc_hd__inv_2 _3803_ (.A(out_data_flat[142]),
    .Y(_1529_));
 sky130_fd_sc_hd__inv_2 _3804_ (.A(out_data_flat[141]),
    .Y(_1530_));
 sky130_fd_sc_hd__inv_2 _3805_ (.A(out_data_flat[140]),
    .Y(_1531_));
 sky130_fd_sc_hd__inv_2 _3806_ (.A(out_data_flat[139]),
    .Y(_1532_));
 sky130_fd_sc_hd__inv_2 _3807_ (.A(out_data_flat[138]),
    .Y(_1533_));
 sky130_fd_sc_hd__inv_2 _3808_ (.A(out_data_flat[137]),
    .Y(_1534_));
 sky130_fd_sc_hd__inv_2 _3809_ (.A(out_data_flat[136]),
    .Y(_1535_));
 sky130_fd_sc_hd__inv_2 _3810_ (.A(out_data_flat[135]),
    .Y(_1536_));
 sky130_fd_sc_hd__inv_2 _3811_ (.A(out_data_flat[134]),
    .Y(_1537_));
 sky130_fd_sc_hd__inv_2 _3812_ (.A(out_data_flat[132]),
    .Y(_1538_));
 sky130_fd_sc_hd__inv_2 _3813_ (.A(out_data_flat[131]),
    .Y(_1539_));
 sky130_fd_sc_hd__inv_2 _3814_ (.A(out_data_flat[130]),
    .Y(_1540_));
 sky130_fd_sc_hd__inv_2 _3815_ (.A(out_data_flat[129]),
    .Y(_1541_));
 sky130_fd_sc_hd__inv_2 _3816_ (.A(out_data_flat[128]),
    .Y(_1542_));
 sky130_fd_sc_hd__inv_2 _3817_ (.A(rst),
    .Y(_0641_));
 sky130_fd_sc_hd__nor2_2 _3818_ (.A(load),
    .B(\gen_pe[1].pe_inst.sel ),
    .Y(_0192_));
 sky130_fd_sc_hd__nor2_2 _3819_ (.A(load),
    .B(_1428_),
    .Y(_1543_));
 sky130_fd_sc_hd__a22o_2 _3820_ (.A1(load),
    .A2(in_data_flat[31]),
    .B1(_0192_),
    .B2(\gen_left[0][31] ),
    .X(_1544_));
 sky130_fd_sc_hd__a21o_2 _3821_ (.A1(out_data_flat[31]),
    .A2(_1543_),
    .B1(_1544_),
    .X(_1409_));
 sky130_fd_sc_hd__a22o_2 _3822_ (.A1(load),
    .A2(in_data_flat[30]),
    .B1(_0192_),
    .B2(\gen_left[0][30] ),
    .X(_1545_));
 sky130_fd_sc_hd__a21o_2 _3823_ (.A1(out_data_flat[30]),
    .A2(_1543_),
    .B1(_1545_),
    .X(_1408_));
 sky130_fd_sc_hd__a22o_2 _3824_ (.A1(load),
    .A2(in_data_flat[29]),
    .B1(_0192_),
    .B2(\gen_left[0][29] ),
    .X(_1546_));
 sky130_fd_sc_hd__a21o_2 _3825_ (.A1(out_data_flat[29]),
    .A2(_1543_),
    .B1(_1546_),
    .X(_1407_));
 sky130_fd_sc_hd__a22o_2 _3826_ (.A1(load),
    .A2(in_data_flat[28]),
    .B1(_0192_),
    .B2(\gen_left[0][28] ),
    .X(_1547_));
 sky130_fd_sc_hd__a21o_2 _3827_ (.A1(out_data_flat[28]),
    .A2(_1543_),
    .B1(_1547_),
    .X(_1406_));
 sky130_fd_sc_hd__a22o_2 _3828_ (.A1(load),
    .A2(in_data_flat[27]),
    .B1(_0192_),
    .B2(\gen_left[0][27] ),
    .X(_1548_));
 sky130_fd_sc_hd__a21o_2 _3829_ (.A1(out_data_flat[27]),
    .A2(_1543_),
    .B1(_1548_),
    .X(_1405_));
 sky130_fd_sc_hd__a22o_2 _3830_ (.A1(load),
    .A2(in_data_flat[26]),
    .B1(_0192_),
    .B2(\gen_left[0][26] ),
    .X(_1549_));
 sky130_fd_sc_hd__a21o_2 _3831_ (.A1(out_data_flat[26]),
    .A2(_1543_),
    .B1(_1549_),
    .X(_1404_));
 sky130_fd_sc_hd__a22o_2 _3832_ (.A1(load),
    .A2(in_data_flat[25]),
    .B1(_0192_),
    .B2(\gen_left[0][25] ),
    .X(_1550_));
 sky130_fd_sc_hd__a21o_2 _3833_ (.A1(out_data_flat[25]),
    .A2(_1543_),
    .B1(_1550_),
    .X(_1403_));
 sky130_fd_sc_hd__a22o_2 _3834_ (.A1(load),
    .A2(in_data_flat[24]),
    .B1(_0192_),
    .B2(\gen_left[0][24] ),
    .X(_1551_));
 sky130_fd_sc_hd__a21o_2 _3835_ (.A1(out_data_flat[24]),
    .A2(_1543_),
    .B1(_1551_),
    .X(_1402_));
 sky130_fd_sc_hd__a22o_2 _3836_ (.A1(load),
    .A2(in_data_flat[23]),
    .B1(_0192_),
    .B2(\gen_left[0][23] ),
    .X(_1552_));
 sky130_fd_sc_hd__a21o_2 _3837_ (.A1(out_data_flat[23]),
    .A2(_1543_),
    .B1(_1552_),
    .X(_1401_));
 sky130_fd_sc_hd__a22o_2 _3838_ (.A1(load),
    .A2(in_data_flat[22]),
    .B1(_0192_),
    .B2(\gen_left[0][22] ),
    .X(_1553_));
 sky130_fd_sc_hd__a21o_2 _3839_ (.A1(out_data_flat[22]),
    .A2(_1543_),
    .B1(_1553_),
    .X(_1400_));
 sky130_fd_sc_hd__a22o_2 _3840_ (.A1(load),
    .A2(in_data_flat[21]),
    .B1(_0192_),
    .B2(\gen_left[0][21] ),
    .X(_1554_));
 sky130_fd_sc_hd__a21o_2 _3841_ (.A1(out_data_flat[21]),
    .A2(_1543_),
    .B1(_1554_),
    .X(_1399_));
 sky130_fd_sc_hd__a22o_2 _3842_ (.A1(load),
    .A2(in_data_flat[20]),
    .B1(_0192_),
    .B2(\gen_left[0][20] ),
    .X(_1555_));
 sky130_fd_sc_hd__a21o_2 _3843_ (.A1(out_data_flat[20]),
    .A2(_1543_),
    .B1(_1555_),
    .X(_1398_));
 sky130_fd_sc_hd__a22o_2 _3844_ (.A1(load),
    .A2(in_data_flat[19]),
    .B1(_0192_),
    .B2(\gen_left[0][19] ),
    .X(_1556_));
 sky130_fd_sc_hd__a21o_2 _3845_ (.A1(out_data_flat[19]),
    .A2(_1543_),
    .B1(_1556_),
    .X(_1397_));
 sky130_fd_sc_hd__a22o_2 _3846_ (.A1(load),
    .A2(in_data_flat[18]),
    .B1(_0192_),
    .B2(\gen_left[0][18] ),
    .X(_1557_));
 sky130_fd_sc_hd__a21o_2 _3847_ (.A1(out_data_flat[18]),
    .A2(_1543_),
    .B1(_1557_),
    .X(_1396_));
 sky130_fd_sc_hd__a22o_2 _3848_ (.A1(load),
    .A2(in_data_flat[17]),
    .B1(_0192_),
    .B2(\gen_left[0][17] ),
    .X(_1558_));
 sky130_fd_sc_hd__a21o_2 _3849_ (.A1(out_data_flat[17]),
    .A2(_1543_),
    .B1(_1558_),
    .X(_1395_));
 sky130_fd_sc_hd__a22o_2 _3850_ (.A1(load),
    .A2(in_data_flat[16]),
    .B1(_0192_),
    .B2(\gen_left[0][16] ),
    .X(_1559_));
 sky130_fd_sc_hd__a21o_2 _3851_ (.A1(out_data_flat[16]),
    .A2(_1543_),
    .B1(_1559_),
    .X(_1394_));
 sky130_fd_sc_hd__a22o_2 _3852_ (.A1(load),
    .A2(in_data_flat[15]),
    .B1(_0192_),
    .B2(\gen_left[0][15] ),
    .X(_1560_));
 sky130_fd_sc_hd__a21o_2 _3853_ (.A1(out_data_flat[15]),
    .A2(_1543_),
    .B1(_1560_),
    .X(_1393_));
 sky130_fd_sc_hd__a22o_2 _3854_ (.A1(load),
    .A2(in_data_flat[14]),
    .B1(_0192_),
    .B2(\gen_left[0][14] ),
    .X(_1561_));
 sky130_fd_sc_hd__a21o_2 _3855_ (.A1(out_data_flat[14]),
    .A2(_1543_),
    .B1(_1561_),
    .X(_1392_));
 sky130_fd_sc_hd__a22o_2 _3856_ (.A1(load),
    .A2(in_data_flat[13]),
    .B1(_0192_),
    .B2(\gen_left[0][13] ),
    .X(_1562_));
 sky130_fd_sc_hd__a21o_2 _3857_ (.A1(out_data_flat[13]),
    .A2(_1543_),
    .B1(_1562_),
    .X(_1391_));
 sky130_fd_sc_hd__a22o_2 _3858_ (.A1(load),
    .A2(in_data_flat[12]),
    .B1(_0192_),
    .B2(\gen_left[0][12] ),
    .X(_1563_));
 sky130_fd_sc_hd__a21o_2 _3859_ (.A1(out_data_flat[12]),
    .A2(_1543_),
    .B1(_1563_),
    .X(_1390_));
 sky130_fd_sc_hd__a22o_2 _3860_ (.A1(load),
    .A2(in_data_flat[11]),
    .B1(_0192_),
    .B2(\gen_left[0][11] ),
    .X(_1564_));
 sky130_fd_sc_hd__a21o_2 _3861_ (.A1(out_data_flat[11]),
    .A2(_1543_),
    .B1(_1564_),
    .X(_1389_));
 sky130_fd_sc_hd__a22o_2 _3862_ (.A1(load),
    .A2(in_data_flat[10]),
    .B1(_0192_),
    .B2(\gen_left[0][10] ),
    .X(_1565_));
 sky130_fd_sc_hd__a21o_2 _3863_ (.A1(out_data_flat[10]),
    .A2(_1543_),
    .B1(_1565_),
    .X(_1388_));
 sky130_fd_sc_hd__a22o_2 _3864_ (.A1(load),
    .A2(in_data_flat[9]),
    .B1(_0192_),
    .B2(\gen_left[0][9] ),
    .X(_1566_));
 sky130_fd_sc_hd__a21o_2 _3865_ (.A1(out_data_flat[9]),
    .A2(_1543_),
    .B1(_1566_),
    .X(_1387_));
 sky130_fd_sc_hd__a22o_2 _3866_ (.A1(load),
    .A2(in_data_flat[8]),
    .B1(_0192_),
    .B2(\gen_left[0][8] ),
    .X(_1567_));
 sky130_fd_sc_hd__a21o_2 _3867_ (.A1(out_data_flat[8]),
    .A2(_1543_),
    .B1(_1567_),
    .X(_1386_));
 sky130_fd_sc_hd__a22o_2 _3868_ (.A1(load),
    .A2(in_data_flat[7]),
    .B1(_0192_),
    .B2(\gen_left[0][7] ),
    .X(_1568_));
 sky130_fd_sc_hd__a21o_2 _3869_ (.A1(out_data_flat[7]),
    .A2(_1543_),
    .B1(_1568_),
    .X(_1385_));
 sky130_fd_sc_hd__a22o_2 _3870_ (.A1(load),
    .A2(in_data_flat[6]),
    .B1(_0192_),
    .B2(\gen_left[0][6] ),
    .X(_1569_));
 sky130_fd_sc_hd__a21o_2 _3871_ (.A1(out_data_flat[6]),
    .A2(_1543_),
    .B1(_1569_),
    .X(_1384_));
 sky130_fd_sc_hd__a22o_2 _3872_ (.A1(load),
    .A2(in_data_flat[5]),
    .B1(_0192_),
    .B2(\gen_left[0][5] ),
    .X(_1570_));
 sky130_fd_sc_hd__a21o_2 _3873_ (.A1(out_data_flat[5]),
    .A2(_1543_),
    .B1(_1570_),
    .X(_1383_));
 sky130_fd_sc_hd__a22o_2 _3874_ (.A1(load),
    .A2(in_data_flat[4]),
    .B1(_0192_),
    .B2(\gen_left[0][4] ),
    .X(_1571_));
 sky130_fd_sc_hd__a21o_2 _3875_ (.A1(out_data_flat[4]),
    .A2(_1543_),
    .B1(_1571_),
    .X(_1382_));
 sky130_fd_sc_hd__a22o_2 _3876_ (.A1(load),
    .A2(in_data_flat[3]),
    .B1(_0192_),
    .B2(\gen_left[0][3] ),
    .X(_1572_));
 sky130_fd_sc_hd__a21o_2 _3877_ (.A1(out_data_flat[3]),
    .A2(_1543_),
    .B1(_1572_),
    .X(_1381_));
 sky130_fd_sc_hd__a22o_2 _3878_ (.A1(load),
    .A2(in_data_flat[2]),
    .B1(_0192_),
    .B2(\gen_left[0][2] ),
    .X(_1573_));
 sky130_fd_sc_hd__a21o_2 _3879_ (.A1(out_data_flat[2]),
    .A2(_1543_),
    .B1(_1573_),
    .X(_1380_));
 sky130_fd_sc_hd__a22o_2 _3880_ (.A1(load),
    .A2(in_data_flat[1]),
    .B1(_0192_),
    .B2(\gen_left[0][1] ),
    .X(_1574_));
 sky130_fd_sc_hd__a21o_2 _3881_ (.A1(out_data_flat[1]),
    .A2(_1543_),
    .B1(_1574_),
    .X(_1379_));
 sky130_fd_sc_hd__a22o_2 _3882_ (.A1(load),
    .A2(in_data_flat[0]),
    .B1(_0192_),
    .B2(\gen_left[0][0] ),
    .X(_1575_));
 sky130_fd_sc_hd__a21o_2 _3883_ (.A1(out_data_flat[0]),
    .A2(_1543_),
    .B1(_1575_),
    .X(_1378_));
 sky130_fd_sc_hd__a22o_2 _3884_ (.A1(load),
    .A2(in_data_flat[255]),
    .B1(_0192_),
    .B2(\gen_pe[6].pe_inst.out_right[31] ),
    .X(_1576_));
 sky130_fd_sc_hd__a21o_2 _3885_ (.A1(out_data_flat[255]),
    .A2(_1543_),
    .B1(_1576_),
    .X(_1377_));
 sky130_fd_sc_hd__a22o_2 _3886_ (.A1(load),
    .A2(in_data_flat[254]),
    .B1(_0192_),
    .B2(\gen_pe[6].pe_inst.out_right[30] ),
    .X(_1577_));
 sky130_fd_sc_hd__a21o_2 _3887_ (.A1(out_data_flat[254]),
    .A2(_1543_),
    .B1(_1577_),
    .X(_1376_));
 sky130_fd_sc_hd__a22o_2 _3888_ (.A1(load),
    .A2(in_data_flat[253]),
    .B1(_0192_),
    .B2(\gen_pe[6].pe_inst.out_right[29] ),
    .X(_1578_));
 sky130_fd_sc_hd__a21o_2 _3889_ (.A1(out_data_flat[253]),
    .A2(_1543_),
    .B1(_1578_),
    .X(_1375_));
 sky130_fd_sc_hd__a22o_2 _3890_ (.A1(load),
    .A2(in_data_flat[252]),
    .B1(_0192_),
    .B2(\gen_pe[6].pe_inst.out_right[28] ),
    .X(_1579_));
 sky130_fd_sc_hd__a21o_2 _3891_ (.A1(out_data_flat[252]),
    .A2(_1543_),
    .B1(_1579_),
    .X(_1374_));
 sky130_fd_sc_hd__a22o_2 _3892_ (.A1(load),
    .A2(in_data_flat[251]),
    .B1(_0192_),
    .B2(\gen_pe[6].pe_inst.out_right[27] ),
    .X(_1580_));
 sky130_fd_sc_hd__a21o_2 _3893_ (.A1(out_data_flat[251]),
    .A2(_1543_),
    .B1(_1580_),
    .X(_1373_));
 sky130_fd_sc_hd__a22o_2 _3894_ (.A1(load),
    .A2(in_data_flat[250]),
    .B1(_0192_),
    .B2(\gen_pe[6].pe_inst.out_right[26] ),
    .X(_1581_));
 sky130_fd_sc_hd__a21o_2 _3895_ (.A1(out_data_flat[250]),
    .A2(_1543_),
    .B1(_1581_),
    .X(_1372_));
 sky130_fd_sc_hd__a22o_2 _3896_ (.A1(load),
    .A2(in_data_flat[249]),
    .B1(_0192_),
    .B2(\gen_pe[6].pe_inst.out_right[25] ),
    .X(_1582_));
 sky130_fd_sc_hd__a21o_2 _3897_ (.A1(out_data_flat[249]),
    .A2(_1543_),
    .B1(_1582_),
    .X(_1371_));
 sky130_fd_sc_hd__a22o_2 _3898_ (.A1(load),
    .A2(in_data_flat[248]),
    .B1(_0192_),
    .B2(\gen_pe[6].pe_inst.out_right[24] ),
    .X(_1583_));
 sky130_fd_sc_hd__a21o_2 _3899_ (.A1(out_data_flat[248]),
    .A2(_1543_),
    .B1(_1583_),
    .X(_1370_));
 sky130_fd_sc_hd__a22o_2 _3900_ (.A1(load),
    .A2(in_data_flat[247]),
    .B1(_0192_),
    .B2(\gen_pe[6].pe_inst.out_right[23] ),
    .X(_1584_));
 sky130_fd_sc_hd__a21o_2 _3901_ (.A1(out_data_flat[247]),
    .A2(_1543_),
    .B1(_1584_),
    .X(_1369_));
 sky130_fd_sc_hd__a22o_2 _3902_ (.A1(load),
    .A2(in_data_flat[246]),
    .B1(_0192_),
    .B2(\gen_pe[6].pe_inst.out_right[22] ),
    .X(_1585_));
 sky130_fd_sc_hd__a21o_2 _3903_ (.A1(out_data_flat[246]),
    .A2(_1543_),
    .B1(_1585_),
    .X(_1368_));
 sky130_fd_sc_hd__a22o_2 _3904_ (.A1(load),
    .A2(in_data_flat[245]),
    .B1(_0192_),
    .B2(\gen_pe[6].pe_inst.out_right[21] ),
    .X(_1586_));
 sky130_fd_sc_hd__a21o_2 _3905_ (.A1(out_data_flat[245]),
    .A2(_1543_),
    .B1(_1586_),
    .X(_1367_));
 sky130_fd_sc_hd__a22o_2 _3906_ (.A1(load),
    .A2(in_data_flat[244]),
    .B1(_0192_),
    .B2(\gen_pe[6].pe_inst.out_right[20] ),
    .X(_1587_));
 sky130_fd_sc_hd__a21o_2 _3907_ (.A1(out_data_flat[244]),
    .A2(_1543_),
    .B1(_1587_),
    .X(_1366_));
 sky130_fd_sc_hd__a22o_2 _3908_ (.A1(load),
    .A2(in_data_flat[243]),
    .B1(_0192_),
    .B2(\gen_pe[6].pe_inst.out_right[19] ),
    .X(_1588_));
 sky130_fd_sc_hd__a21o_2 _3909_ (.A1(out_data_flat[243]),
    .A2(_1543_),
    .B1(_1588_),
    .X(_1365_));
 sky130_fd_sc_hd__a22o_2 _3910_ (.A1(load),
    .A2(in_data_flat[242]),
    .B1(_0192_),
    .B2(\gen_pe[6].pe_inst.out_right[18] ),
    .X(_1589_));
 sky130_fd_sc_hd__a21o_2 _3911_ (.A1(out_data_flat[242]),
    .A2(_1543_),
    .B1(_1589_),
    .X(_1364_));
 sky130_fd_sc_hd__a22o_2 _3912_ (.A1(load),
    .A2(in_data_flat[241]),
    .B1(_0192_),
    .B2(\gen_pe[6].pe_inst.out_right[17] ),
    .X(_1590_));
 sky130_fd_sc_hd__a21o_2 _3913_ (.A1(out_data_flat[241]),
    .A2(_1543_),
    .B1(_1590_),
    .X(_1363_));
 sky130_fd_sc_hd__a22o_2 _3914_ (.A1(load),
    .A2(in_data_flat[240]),
    .B1(_0192_),
    .B2(\gen_pe[6].pe_inst.out_right[16] ),
    .X(_1591_));
 sky130_fd_sc_hd__a21o_2 _3915_ (.A1(out_data_flat[240]),
    .A2(_1543_),
    .B1(_1591_),
    .X(_1362_));
 sky130_fd_sc_hd__a22o_2 _3916_ (.A1(load),
    .A2(in_data_flat[239]),
    .B1(_0192_),
    .B2(\gen_pe[6].pe_inst.out_right[15] ),
    .X(_1592_));
 sky130_fd_sc_hd__a21o_2 _3917_ (.A1(out_data_flat[239]),
    .A2(_1543_),
    .B1(_1592_),
    .X(_1361_));
 sky130_fd_sc_hd__a22o_2 _3918_ (.A1(load),
    .A2(in_data_flat[238]),
    .B1(_0192_),
    .B2(\gen_pe[6].pe_inst.out_right[14] ),
    .X(_1593_));
 sky130_fd_sc_hd__a21o_2 _3919_ (.A1(out_data_flat[238]),
    .A2(_1543_),
    .B1(_1593_),
    .X(_1360_));
 sky130_fd_sc_hd__a22o_2 _3920_ (.A1(load),
    .A2(in_data_flat[237]),
    .B1(_0192_),
    .B2(\gen_pe[6].pe_inst.out_right[13] ),
    .X(_1594_));
 sky130_fd_sc_hd__a21o_2 _3921_ (.A1(out_data_flat[237]),
    .A2(_1543_),
    .B1(_1594_),
    .X(_1359_));
 sky130_fd_sc_hd__a22o_2 _3922_ (.A1(load),
    .A2(in_data_flat[236]),
    .B1(_0192_),
    .B2(\gen_pe[6].pe_inst.out_right[12] ),
    .X(_1595_));
 sky130_fd_sc_hd__a21o_2 _3923_ (.A1(out_data_flat[236]),
    .A2(_1543_),
    .B1(_1595_),
    .X(_1358_));
 sky130_fd_sc_hd__a22o_2 _3924_ (.A1(load),
    .A2(in_data_flat[235]),
    .B1(_0192_),
    .B2(\gen_pe[6].pe_inst.out_right[11] ),
    .X(_1596_));
 sky130_fd_sc_hd__a21o_2 _3925_ (.A1(out_data_flat[235]),
    .A2(_1543_),
    .B1(_1596_),
    .X(_1357_));
 sky130_fd_sc_hd__a22o_2 _3926_ (.A1(load),
    .A2(in_data_flat[234]),
    .B1(_0192_),
    .B2(\gen_pe[6].pe_inst.out_right[10] ),
    .X(_1597_));
 sky130_fd_sc_hd__a21o_2 _3927_ (.A1(out_data_flat[234]),
    .A2(_1543_),
    .B1(_1597_),
    .X(_1356_));
 sky130_fd_sc_hd__a22o_2 _3928_ (.A1(load),
    .A2(in_data_flat[233]),
    .B1(_0192_),
    .B2(\gen_pe[6].pe_inst.out_right[9] ),
    .X(_1598_));
 sky130_fd_sc_hd__a21o_2 _3929_ (.A1(out_data_flat[233]),
    .A2(_1543_),
    .B1(_1598_),
    .X(_1355_));
 sky130_fd_sc_hd__a22o_2 _3930_ (.A1(load),
    .A2(in_data_flat[232]),
    .B1(_0192_),
    .B2(\gen_pe[6].pe_inst.out_right[8] ),
    .X(_1599_));
 sky130_fd_sc_hd__a21o_2 _3931_ (.A1(out_data_flat[232]),
    .A2(_1543_),
    .B1(_1599_),
    .X(_1354_));
 sky130_fd_sc_hd__a22o_2 _3932_ (.A1(load),
    .A2(in_data_flat[231]),
    .B1(_0192_),
    .B2(\gen_pe[6].pe_inst.out_right[7] ),
    .X(_1600_));
 sky130_fd_sc_hd__a21o_2 _3933_ (.A1(out_data_flat[231]),
    .A2(_1543_),
    .B1(_1600_),
    .X(_1353_));
 sky130_fd_sc_hd__a22o_2 _3934_ (.A1(load),
    .A2(in_data_flat[230]),
    .B1(_0192_),
    .B2(\gen_pe[6].pe_inst.out_right[6] ),
    .X(_1601_));
 sky130_fd_sc_hd__a21o_2 _3935_ (.A1(out_data_flat[230]),
    .A2(_1543_),
    .B1(_1601_),
    .X(_1352_));
 sky130_fd_sc_hd__a22o_2 _3936_ (.A1(load),
    .A2(in_data_flat[229]),
    .B1(_0192_),
    .B2(\gen_pe[6].pe_inst.out_right[5] ),
    .X(_1602_));
 sky130_fd_sc_hd__a21o_2 _3937_ (.A1(out_data_flat[229]),
    .A2(_1543_),
    .B1(_1602_),
    .X(_1351_));
 sky130_fd_sc_hd__a22o_2 _3938_ (.A1(load),
    .A2(in_data_flat[228]),
    .B1(_0192_),
    .B2(\gen_pe[6].pe_inst.out_right[4] ),
    .X(_1603_));
 sky130_fd_sc_hd__a21o_2 _3939_ (.A1(out_data_flat[228]),
    .A2(_1543_),
    .B1(_1603_),
    .X(_1350_));
 sky130_fd_sc_hd__a22o_2 _3940_ (.A1(load),
    .A2(in_data_flat[227]),
    .B1(_0192_),
    .B2(\gen_pe[6].pe_inst.out_right[3] ),
    .X(_1604_));
 sky130_fd_sc_hd__a21o_2 _3941_ (.A1(out_data_flat[227]),
    .A2(_1543_),
    .B1(_1604_),
    .X(_1349_));
 sky130_fd_sc_hd__a22o_2 _3942_ (.A1(load),
    .A2(in_data_flat[226]),
    .B1(_0192_),
    .B2(\gen_pe[6].pe_inst.out_right[2] ),
    .X(_1605_));
 sky130_fd_sc_hd__a21o_2 _3943_ (.A1(out_data_flat[226]),
    .A2(_1543_),
    .B1(_1605_),
    .X(_1348_));
 sky130_fd_sc_hd__a22o_2 _3944_ (.A1(load),
    .A2(in_data_flat[225]),
    .B1(_0192_),
    .B2(\gen_pe[6].pe_inst.out_right[1] ),
    .X(_1606_));
 sky130_fd_sc_hd__a21o_2 _3945_ (.A1(out_data_flat[225]),
    .A2(_1543_),
    .B1(_1606_),
    .X(_1347_));
 sky130_fd_sc_hd__a22o_2 _3946_ (.A1(load),
    .A2(in_data_flat[224]),
    .B1(_0192_),
    .B2(\gen_pe[6].pe_inst.out_right[0] ),
    .X(_1607_));
 sky130_fd_sc_hd__a21o_2 _3947_ (.A1(out_data_flat[224]),
    .A2(_1543_),
    .B1(_1607_),
    .X(_1346_));
 sky130_fd_sc_hd__a22o_2 _3948_ (.A1(out_data_flat[29]),
    .A2(_1431_),
    .B1(_1432_),
    .B2(out_data_flat[28]),
    .X(_1608_));
 sky130_fd_sc_hd__and2b_2 _3949_ (.A_N(out_data_flat[31]),
    .B(out_data_flat[63]),
    .X(_1609_));
 sky130_fd_sc_hd__o21bai_2 _3950_ (.A1(out_data_flat[28]),
    .A2(_1432_),
    .B1_N(_1609_),
    .Y(_1610_));
 sky130_fd_sc_hd__a22o_2 _3951_ (.A1(out_data_flat[31]),
    .A2(_1429_),
    .B1(_1430_),
    .B2(out_data_flat[30]),
    .X(_1611_));
 sky130_fd_sc_hd__o22a_2 _3952_ (.A1(out_data_flat[30]),
    .A2(_1430_),
    .B1(_1431_),
    .B2(out_data_flat[29]),
    .X(_1612_));
 sky130_fd_sc_hd__or4b_2 _3953_ (.A(_1608_),
    .B(_1610_),
    .C(_1611_),
    .D_N(_1612_),
    .X(_1613_));
 sky130_fd_sc_hd__xor2_2 _3954_ (.A(out_data_flat[26]),
    .B(out_data_flat[58]),
    .X(_1614_));
 sky130_fd_sc_hd__and2b_2 _3955_ (.A_N(out_data_flat[27]),
    .B(out_data_flat[59]),
    .X(_1615_));
 sky130_fd_sc_hd__nand2b_2 _3956_ (.A_N(out_data_flat[59]),
    .B(out_data_flat[27]),
    .Y(_1616_));
 sky130_fd_sc_hd__nor2_2 _3957_ (.A(out_data_flat[25]),
    .B(_1433_),
    .Y(_1617_));
 sky130_fd_sc_hd__or3b_2 _3958_ (.A(_1614_),
    .B(_1615_),
    .C_N(_1616_),
    .X(_1618_));
 sky130_fd_sc_hd__a2bb2o_2 _3959_ (.A1_N(out_data_flat[56]),
    .A2_N(_1411_),
    .B1(out_data_flat[25]),
    .B2(_1433_),
    .X(_1619_));
 sky130_fd_sc_hd__a2111o_2 _3960_ (.A1(_1411_),
    .A2(out_data_flat[56]),
    .B1(_1617_),
    .C1(_1618_),
    .D1(_1619_),
    .X(_1620_));
 sky130_fd_sc_hd__nor2_2 _3961_ (.A(_1613_),
    .B(_1620_),
    .Y(_1621_));
 sky130_fd_sc_hd__a22o_2 _3962_ (.A1(out_data_flat[19]),
    .A2(_1438_),
    .B1(_1439_),
    .B2(out_data_flat[18]),
    .X(_1622_));
 sky130_fd_sc_hd__nand2b_2 _3963_ (.A_N(out_data_flat[19]),
    .B(out_data_flat[51]),
    .Y(_1623_));
 sky130_fd_sc_hd__o221a_2 _3964_ (.A1(out_data_flat[18]),
    .A2(_1439_),
    .B1(_1440_),
    .B2(out_data_flat[17]),
    .C1(_1623_),
    .X(_1624_));
 sky130_fd_sc_hd__and2b_2 _3965_ (.A_N(_1622_),
    .B(_1624_),
    .X(_1625_));
 sky130_fd_sc_hd__a22o_2 _3966_ (.A1(out_data_flat[23]),
    .A2(_1434_),
    .B1(_1435_),
    .B2(out_data_flat[22]),
    .X(_1626_));
 sky130_fd_sc_hd__a22o_2 _3967_ (.A1(out_data_flat[21]),
    .A2(_1436_),
    .B1(_1437_),
    .B2(out_data_flat[20]),
    .X(_1627_));
 sky130_fd_sc_hd__nor2_2 _3968_ (.A(out_data_flat[23]),
    .B(_1434_),
    .Y(_1628_));
 sky130_fd_sc_hd__o21ba_2 _3969_ (.A1(out_data_flat[20]),
    .A2(_1437_),
    .B1_N(_1628_),
    .X(_1629_));
 sky130_fd_sc_hd__o22a_2 _3970_ (.A1(out_data_flat[22]),
    .A2(_1435_),
    .B1(_1436_),
    .B2(out_data_flat[21]),
    .X(_1630_));
 sky130_fd_sc_hd__and4bb_2 _3971_ (.A_N(_1626_),
    .B_N(_1627_),
    .C(_1629_),
    .D(_1630_),
    .X(_1631_));
 sky130_fd_sc_hd__a22o_2 _3972_ (.A1(out_data_flat[17]),
    .A2(_1440_),
    .B1(_1441_),
    .B2(out_data_flat[16]),
    .X(_1632_));
 sky130_fd_sc_hd__o21ba_2 _3973_ (.A1(out_data_flat[16]),
    .A2(_1441_),
    .B1_N(_1632_),
    .X(_1633_));
 sky130_fd_sc_hd__nand4_2 _3974_ (.A(_1621_),
    .B(_1625_),
    .C(_1631_),
    .D(_1633_),
    .Y(_1634_));
 sky130_fd_sc_hd__nand2b_2 _3975_ (.A_N(out_data_flat[47]),
    .B(out_data_flat[15]),
    .Y(_1635_));
 sky130_fd_sc_hd__o21ai_2 _3976_ (.A1(_1412_),
    .A2(out_data_flat[46]),
    .B1(_1635_),
    .Y(_1636_));
 sky130_fd_sc_hd__nand2b_2 _3977_ (.A_N(out_data_flat[15]),
    .B(out_data_flat[47]),
    .Y(_1637_));
 sky130_fd_sc_hd__xnor2_2 _3978_ (.A(out_data_flat[14]),
    .B(out_data_flat[46]),
    .Y(_1638_));
 sky130_fd_sc_hd__and3_2 _3979_ (.A(_1635_),
    .B(_1637_),
    .C(_1638_),
    .X(_1639_));
 sky130_fd_sc_hd__a22o_2 _3980_ (.A1(out_data_flat[13]),
    .A2(_1443_),
    .B1(_1444_),
    .B2(out_data_flat[12]),
    .X(_1640_));
 sky130_fd_sc_hd__or2_2 _3981_ (.A(out_data_flat[13]),
    .B(_1443_),
    .X(_1641_));
 sky130_fd_sc_hd__nor2_2 _3982_ (.A(out_data_flat[12]),
    .B(_1444_),
    .Y(_1642_));
 sky130_fd_sc_hd__or4bb_2 _3983_ (.A(_1642_),
    .B(_1640_),
    .C_N(_1639_),
    .D_N(_1641_),
    .X(_1643_));
 sky130_fd_sc_hd__nand2b_2 _3984_ (.A_N(out_data_flat[43]),
    .B(out_data_flat[11]),
    .Y(_1644_));
 sky130_fd_sc_hd__and2b_2 _3985_ (.A_N(out_data_flat[11]),
    .B(out_data_flat[43]),
    .X(_1645_));
 sky130_fd_sc_hd__xor2_2 _3986_ (.A(out_data_flat[10]),
    .B(out_data_flat[42]),
    .X(_1646_));
 sky130_fd_sc_hd__or3b_2 _3987_ (.A(_1646_),
    .B(_1645_),
    .C_N(_1644_),
    .X(_1647_));
 sky130_fd_sc_hd__o22a_2 _3988_ (.A1(_1413_),
    .A2(out_data_flat[41]),
    .B1(out_data_flat[40]),
    .B2(_1414_),
    .X(_1648_));
 sky130_fd_sc_hd__and2_2 _3989_ (.A(_1413_),
    .B(out_data_flat[41]),
    .X(_1649_));
 sky130_fd_sc_hd__and2_2 _3990_ (.A(_1414_),
    .B(out_data_flat[40]),
    .X(_1650_));
 sky130_fd_sc_hd__or4b_2 _3991_ (.A(_1647_),
    .B(_1649_),
    .C(_1650_),
    .D_N(_1648_),
    .X(_1651_));
 sky130_fd_sc_hd__a2bb2o_2 _3992_ (.A1_N(out_data_flat[36]),
    .A2_N(_1415_),
    .B1(out_data_flat[5]),
    .B2(_1447_),
    .X(_1652_));
 sky130_fd_sc_hd__nand2b_2 _3993_ (.A_N(out_data_flat[39]),
    .B(out_data_flat[7]),
    .Y(_1653_));
 sky130_fd_sc_hd__nor2_2 _3994_ (.A(out_data_flat[5]),
    .B(_1447_),
    .Y(_1654_));
 sky130_fd_sc_hd__and2b_2 _3995_ (.A_N(out_data_flat[7]),
    .B(out_data_flat[39]),
    .X(_1655_));
 sky130_fd_sc_hd__xor2_2 _3996_ (.A(out_data_flat[6]),
    .B(out_data_flat[38]),
    .X(_1656_));
 sky130_fd_sc_hd__or3b_2 _3997_ (.A(_1656_),
    .B(_1655_),
    .C_N(_1653_),
    .X(_1657_));
 sky130_fd_sc_hd__or3b_2 _3998_ (.A(_1657_),
    .B(_1654_),
    .C_N(_1652_),
    .X(_1658_));
 sky130_fd_sc_hd__or3b_2 _3999_ (.A(out_data_flat[38]),
    .B(_1655_),
    .C_N(out_data_flat[6]),
    .X(_1659_));
 sky130_fd_sc_hd__a311o_2 _4000_ (.A1(_1653_),
    .A2(_1658_),
    .A3(_1659_),
    .B1(_1651_),
    .C1(_1643_),
    .X(_1660_));
 sky130_fd_sc_hd__a2111o_2 _4001_ (.A1(_1415_),
    .A2(out_data_flat[36]),
    .B1(_1652_),
    .C1(_1654_),
    .D1(_1657_),
    .X(_1661_));
 sky130_fd_sc_hd__or3_2 _4002_ (.A(_1643_),
    .B(_1651_),
    .C(_1661_),
    .X(_1662_));
 sky130_fd_sc_hd__and2b_2 _4003_ (.A_N(out_data_flat[3]),
    .B(out_data_flat[35]),
    .X(_1663_));
 sky130_fd_sc_hd__nand2b_2 _4004_ (.A_N(out_data_flat[35]),
    .B(out_data_flat[3]),
    .Y(_1664_));
 sky130_fd_sc_hd__o21ai_2 _4005_ (.A1(out_data_flat[2]),
    .A2(_1448_),
    .B1(_1664_),
    .Y(_1665_));
 sky130_fd_sc_hd__a211o_2 _4006_ (.A1(out_data_flat[2]),
    .A2(_1448_),
    .B1(_1663_),
    .C1(_1665_),
    .X(_1666_));
 sky130_fd_sc_hd__or2_2 _4007_ (.A(_1416_),
    .B(out_data_flat[33]),
    .X(_1667_));
 sky130_fd_sc_hd__a22o_2 _4008_ (.A1(_1416_),
    .A2(out_data_flat[33]),
    .B1(out_data_flat[32]),
    .B2(_1417_),
    .X(_1668_));
 sky130_fd_sc_hd__a21o_2 _4009_ (.A1(_1667_),
    .A2(_1668_),
    .B1(_1666_),
    .X(_1669_));
 sky130_fd_sc_hd__or3b_2 _4010_ (.A(out_data_flat[34]),
    .B(_1663_),
    .C_N(out_data_flat[2]),
    .X(_1670_));
 sky130_fd_sc_hd__a31o_2 _4011_ (.A1(_1664_),
    .A2(_1669_),
    .A3(_1670_),
    .B1(_1662_),
    .X(_1671_));
 sky130_fd_sc_hd__or3_2 _4012_ (.A(_1647_),
    .B(_1648_),
    .C(_1649_),
    .X(_1672_));
 sky130_fd_sc_hd__or3b_2 _4013_ (.A(out_data_flat[42]),
    .B(_1645_),
    .C_N(out_data_flat[10]),
    .X(_1673_));
 sky130_fd_sc_hd__a31o_2 _4014_ (.A1(_1644_),
    .A2(_1672_),
    .A3(_1673_),
    .B1(_1643_),
    .X(_1674_));
 sky130_fd_sc_hd__a32oi_2 _4015_ (.A1(_1639_),
    .A2(_1640_),
    .A3(_1641_),
    .B1(_1637_),
    .B2(_1636_),
    .Y(_1675_));
 sky130_fd_sc_hd__a41o_2 _4016_ (.A1(_1660_),
    .A2(_1671_),
    .A3(_1674_),
    .A4(_1675_),
    .B1(_1634_),
    .X(_1676_));
 sky130_fd_sc_hd__a21oi_2 _4017_ (.A1(_1627_),
    .A2(_1630_),
    .B1(_1626_),
    .Y(_1677_));
 sky130_fd_sc_hd__o211a_2 _4018_ (.A1(out_data_flat[19]),
    .A2(_1438_),
    .B1(_1439_),
    .C1(out_data_flat[18]),
    .X(_1678_));
 sky130_fd_sc_hd__a221o_2 _4019_ (.A1(out_data_flat[19]),
    .A2(_1438_),
    .B1(_1625_),
    .B2(_1632_),
    .C1(_1678_),
    .X(_1679_));
 sky130_fd_sc_hd__a2bb2o_2 _4020_ (.A1_N(_1628_),
    .A2_N(_1677_),
    .B1(_1679_),
    .B2(_1631_),
    .X(_1680_));
 sky130_fd_sc_hd__nand2_2 _4021_ (.A(_1621_),
    .B(_1680_),
    .Y(_1681_));
 sky130_fd_sc_hd__or4b_2 _4022_ (.A(_1613_),
    .B(_1617_),
    .C(_1618_),
    .D_N(_1619_),
    .X(_1682_));
 sky130_fd_sc_hd__a21oi_2 _4023_ (.A1(_1608_),
    .A2(_1612_),
    .B1(_1611_),
    .Y(_1683_));
 sky130_fd_sc_hd__o31a_2 _4024_ (.A1(_1410_),
    .A2(out_data_flat[58]),
    .A3(_1615_),
    .B1(_1616_),
    .X(_1684_));
 sky130_fd_sc_hd__o221a_2 _4025_ (.A1(_1609_),
    .A2(_1683_),
    .B1(_1684_),
    .B2(_1613_),
    .C1(_1682_),
    .X(_1685_));
 sky130_fd_sc_hd__o21ai_2 _4026_ (.A1(_1417_),
    .A2(out_data_flat[32]),
    .B1(_1667_),
    .Y(_1686_));
 sky130_fd_sc_hd__or4_2 _4027_ (.A(_1662_),
    .B(_1666_),
    .C(_1668_),
    .D(_1686_),
    .X(_1687_));
 sky130_fd_sc_hd__nor2_2 _4028_ (.A(_1634_),
    .B(_1687_),
    .Y(_1688_));
 sky130_fd_sc_hd__a311o_2 _4029_ (.A1(_1676_),
    .A2(_1681_),
    .A3(_1685_),
    .B1(_1688_),
    .C1(\gen_pe[1].pe_inst.sel ),
    .X(_1689_));
 sky130_fd_sc_hd__mux2_1 _4030_ (.A0(out_data_flat[0]),
    .A1(out_data_flat[32]),
    .S(_1689_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _4031_ (.A0(out_data_flat[1]),
    .A1(out_data_flat[33]),
    .S(_1689_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _4032_ (.A0(out_data_flat[2]),
    .A1(out_data_flat[34]),
    .S(_1689_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _4033_ (.A0(out_data_flat[3]),
    .A1(out_data_flat[35]),
    .S(_1689_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _4034_ (.A0(out_data_flat[4]),
    .A1(out_data_flat[36]),
    .S(_1689_),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _4035_ (.A0(out_data_flat[5]),
    .A1(out_data_flat[37]),
    .S(_1689_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _4036_ (.A0(out_data_flat[6]),
    .A1(out_data_flat[38]),
    .S(_1689_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _4037_ (.A0(out_data_flat[7]),
    .A1(out_data_flat[39]),
    .S(_1689_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _4038_ (.A0(out_data_flat[8]),
    .A1(out_data_flat[40]),
    .S(_1689_),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _4039_ (.A0(out_data_flat[9]),
    .A1(out_data_flat[41]),
    .S(_1689_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _4040_ (.A0(out_data_flat[10]),
    .A1(out_data_flat[42]),
    .S(_1689_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _4041_ (.A0(out_data_flat[11]),
    .A1(out_data_flat[43]),
    .S(_1689_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _4042_ (.A0(out_data_flat[12]),
    .A1(out_data_flat[44]),
    .S(_1689_),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _4043_ (.A0(out_data_flat[13]),
    .A1(out_data_flat[45]),
    .S(_1689_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _4044_ (.A0(out_data_flat[14]),
    .A1(out_data_flat[46]),
    .S(_1689_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _4045_ (.A0(out_data_flat[15]),
    .A1(out_data_flat[47]),
    .S(_1689_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _4046_ (.A0(out_data_flat[16]),
    .A1(out_data_flat[48]),
    .S(_1689_),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _4047_ (.A0(out_data_flat[17]),
    .A1(out_data_flat[49]),
    .S(_1689_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _4048_ (.A0(out_data_flat[18]),
    .A1(out_data_flat[50]),
    .S(_1689_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _4049_ (.A0(out_data_flat[19]),
    .A1(out_data_flat[51]),
    .S(_1689_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _4050_ (.A0(out_data_flat[20]),
    .A1(out_data_flat[52]),
    .S(_1689_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _4051_ (.A0(out_data_flat[21]),
    .A1(out_data_flat[53]),
    .S(_1689_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _4052_ (.A0(out_data_flat[22]),
    .A1(out_data_flat[54]),
    .S(_1689_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _4053_ (.A0(out_data_flat[23]),
    .A1(out_data_flat[55]),
    .S(_1689_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _4054_ (.A0(out_data_flat[24]),
    .A1(out_data_flat[56]),
    .S(_1689_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _4055_ (.A0(out_data_flat[25]),
    .A1(out_data_flat[57]),
    .S(_1689_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _4056_ (.A0(out_data_flat[26]),
    .A1(out_data_flat[58]),
    .S(_1689_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _4057_ (.A0(out_data_flat[27]),
    .A1(out_data_flat[59]),
    .S(_1689_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _4058_ (.A0(out_data_flat[28]),
    .A1(out_data_flat[60]),
    .S(_1689_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _4059_ (.A0(out_data_flat[29]),
    .A1(out_data_flat[61]),
    .S(_1689_),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _4060_ (.A0(out_data_flat[30]),
    .A1(out_data_flat[62]),
    .S(_1689_),
    .X(_0248_));
 sky130_fd_sc_hd__a21o_2 _4061_ (.A1(out_data_flat[31]),
    .A2(_1428_),
    .B1(out_data_flat[63]),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _4062_ (.A0(out_data_flat[32]),
    .A1(out_data_flat[0]),
    .S(_1689_),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _4063_ (.A0(out_data_flat[33]),
    .A1(out_data_flat[1]),
    .S(_1689_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _4064_ (.A0(out_data_flat[34]),
    .A1(out_data_flat[2]),
    .S(_1689_),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _4065_ (.A0(out_data_flat[35]),
    .A1(out_data_flat[3]),
    .S(_1689_),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _4066_ (.A0(out_data_flat[36]),
    .A1(out_data_flat[4]),
    .S(_1689_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _4067_ (.A0(out_data_flat[37]),
    .A1(out_data_flat[5]),
    .S(_1689_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _4068_ (.A0(out_data_flat[38]),
    .A1(out_data_flat[6]),
    .S(_1689_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _4069_ (.A0(out_data_flat[39]),
    .A1(out_data_flat[7]),
    .S(_1689_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _4070_ (.A0(out_data_flat[40]),
    .A1(out_data_flat[8]),
    .S(_1689_),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _4071_ (.A0(out_data_flat[41]),
    .A1(out_data_flat[9]),
    .S(_1689_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _4072_ (.A0(out_data_flat[42]),
    .A1(out_data_flat[10]),
    .S(_1689_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _4073_ (.A0(out_data_flat[43]),
    .A1(out_data_flat[11]),
    .S(_1689_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _4074_ (.A0(out_data_flat[44]),
    .A1(out_data_flat[12]),
    .S(_1689_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _4075_ (.A0(out_data_flat[45]),
    .A1(out_data_flat[13]),
    .S(_1689_),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _4076_ (.A0(out_data_flat[46]),
    .A1(out_data_flat[14]),
    .S(_1689_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _4077_ (.A0(out_data_flat[47]),
    .A1(out_data_flat[15]),
    .S(_1689_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _4078_ (.A0(out_data_flat[48]),
    .A1(out_data_flat[16]),
    .S(_1689_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _4079_ (.A0(out_data_flat[49]),
    .A1(out_data_flat[17]),
    .S(_1689_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _4080_ (.A0(out_data_flat[50]),
    .A1(out_data_flat[18]),
    .S(_1689_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _4081_ (.A0(out_data_flat[51]),
    .A1(out_data_flat[19]),
    .S(_1689_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _4082_ (.A0(out_data_flat[52]),
    .A1(out_data_flat[20]),
    .S(_1689_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _4083_ (.A0(out_data_flat[53]),
    .A1(out_data_flat[21]),
    .S(_1689_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _4084_ (.A0(out_data_flat[54]),
    .A1(out_data_flat[22]),
    .S(_1689_),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _4085_ (.A0(out_data_flat[55]),
    .A1(out_data_flat[23]),
    .S(_1689_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _4086_ (.A0(out_data_flat[56]),
    .A1(out_data_flat[24]),
    .S(_1689_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _4087_ (.A0(out_data_flat[57]),
    .A1(out_data_flat[25]),
    .S(_1689_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _4088_ (.A0(out_data_flat[58]),
    .A1(out_data_flat[26]),
    .S(_1689_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _4089_ (.A0(out_data_flat[59]),
    .A1(out_data_flat[27]),
    .S(_1689_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _4090_ (.A0(out_data_flat[60]),
    .A1(out_data_flat[28]),
    .S(_1689_),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _4091_ (.A0(out_data_flat[61]),
    .A1(out_data_flat[29]),
    .S(_1689_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _4092_ (.A0(out_data_flat[62]),
    .A1(out_data_flat[30]),
    .S(_1689_),
    .X(_0216_));
 sky130_fd_sc_hd__o21a_2 _4093_ (.A1(\gen_pe[1].pe_inst.sel ),
    .A2(out_data_flat[63]),
    .B1(out_data_flat[31]),
    .X(_0217_));
 sky130_fd_sc_hd__xor2_2 _4094_ (.A(out_data_flat[255]),
    .B(out_data_flat[223]),
    .X(_1690_));
 sky130_fd_sc_hd__nand2_2 _4095_ (.A(out_data_flat[254]),
    .B(_1450_),
    .Y(_1691_));
 sky130_fd_sc_hd__o22a_2 _4096_ (.A1(out_data_flat[254]),
    .A2(_1450_),
    .B1(_1451_),
    .B2(out_data_flat[253]),
    .X(_1692_));
 sky130_fd_sc_hd__and3b_2 _4097_ (.A_N(_1690_),
    .B(_1691_),
    .C(_1692_),
    .X(_1693_));
 sky130_fd_sc_hd__a22o_2 _4098_ (.A1(out_data_flat[253]),
    .A2(_1451_),
    .B1(_1452_),
    .B2(out_data_flat[252]),
    .X(_1694_));
 sky130_fd_sc_hd__inv_2 _4099_ (.A(_1694_),
    .Y(_1695_));
 sky130_fd_sc_hd__o211a_2 _4100_ (.A1(out_data_flat[252]),
    .A2(_1452_),
    .B1(_1693_),
    .C1(_1695_),
    .X(_1696_));
 sky130_fd_sc_hd__o22a_2 _4101_ (.A1(_1419_),
    .A2(out_data_flat[219]),
    .B1(out_data_flat[218]),
    .B2(_1420_),
    .X(_1697_));
 sky130_fd_sc_hd__and2_2 _4102_ (.A(_1419_),
    .B(out_data_flat[219]),
    .X(_1698_));
 sky130_fd_sc_hd__and2_2 _4103_ (.A(_1420_),
    .B(out_data_flat[218]),
    .X(_1699_));
 sky130_fd_sc_hd__and2_2 _4104_ (.A(_1421_),
    .B(out_data_flat[217]),
    .X(_1700_));
 sky130_fd_sc_hd__or3b_2 _4105_ (.A(_1698_),
    .B(_1699_),
    .C_N(_1697_),
    .X(_1701_));
 sky130_fd_sc_hd__nor2_2 _4106_ (.A(_1700_),
    .B(_1701_),
    .Y(_1702_));
 sky130_fd_sc_hd__o2bb2a_2 _4107_ (.A1_N(_1453_),
    .A2_N(out_data_flat[248]),
    .B1(_1421_),
    .B2(out_data_flat[217]),
    .X(_1703_));
 sky130_fd_sc_hd__o2111a_2 _4108_ (.A1(out_data_flat[248]),
    .A2(_1453_),
    .B1(_1696_),
    .C1(_1702_),
    .D1(_1703_),
    .X(_1704_));
 sky130_fd_sc_hd__o2bb2a_2 _4109_ (.A1_N(_1457_),
    .A2_N(out_data_flat[240]),
    .B1(_1423_),
    .B2(out_data_flat[209]),
    .X(_1705_));
 sky130_fd_sc_hd__and2b_2 _4110_ (.A_N(out_data_flat[215]),
    .B(out_data_flat[247]),
    .X(_1706_));
 sky130_fd_sc_hd__and2b_2 _4111_ (.A_N(out_data_flat[214]),
    .B(out_data_flat[246]),
    .X(_1707_));
 sky130_fd_sc_hd__nor2_2 _4112_ (.A(_1706_),
    .B(_1707_),
    .Y(_1708_));
 sky130_fd_sc_hd__and2b_2 _4113_ (.A_N(out_data_flat[247]),
    .B(out_data_flat[215]),
    .X(_1709_));
 sky130_fd_sc_hd__nor2_2 _4114_ (.A(out_data_flat[245]),
    .B(_1454_),
    .Y(_1710_));
 sky130_fd_sc_hd__and2b_2 _4115_ (.A_N(out_data_flat[246]),
    .B(out_data_flat[214]),
    .X(_1711_));
 sky130_fd_sc_hd__or4_2 _4116_ (.A(_1706_),
    .B(_1707_),
    .C(_1709_),
    .D(_1711_),
    .X(_1712_));
 sky130_fd_sc_hd__o2bb2a_2 _4117_ (.A1_N(out_data_flat[245]),
    .A2_N(_1454_),
    .B1(out_data_flat[212]),
    .B2(_1422_),
    .X(_1713_));
 sky130_fd_sc_hd__nand2_2 _4118_ (.A(_1422_),
    .B(out_data_flat[212]),
    .Y(_1714_));
 sky130_fd_sc_hd__and4bb_2 _4119_ (.A_N(_1710_),
    .B_N(_1712_),
    .C(_1713_),
    .D(_1714_),
    .X(_1715_));
 sky130_fd_sc_hd__nand2b_2 _4120_ (.A_N(out_data_flat[243]),
    .B(out_data_flat[211]),
    .Y(_1716_));
 sky130_fd_sc_hd__and2b_2 _4121_ (.A_N(out_data_flat[241]),
    .B(out_data_flat[209]),
    .X(_1717_));
 sky130_fd_sc_hd__and2b_2 _4122_ (.A_N(out_data_flat[211]),
    .B(out_data_flat[243]),
    .X(_1718_));
 sky130_fd_sc_hd__xor2_2 _4123_ (.A(out_data_flat[242]),
    .B(out_data_flat[210]),
    .X(_1719_));
 sky130_fd_sc_hd__or4b_2 _4124_ (.A(_1717_),
    .B(_1719_),
    .C(_1718_),
    .D_N(_1716_),
    .X(_1720_));
 sky130_fd_sc_hd__inv_2 _4125_ (.A(_1720_),
    .Y(_1721_));
 sky130_fd_sc_hd__a31o_2 _4126_ (.A1(out_data_flat[242]),
    .A2(_1456_),
    .A3(_1716_),
    .B1(_1718_),
    .X(_1722_));
 sky130_fd_sc_hd__or3_2 _4127_ (.A(_1710_),
    .B(_1712_),
    .C(_1713_),
    .X(_1723_));
 sky130_fd_sc_hd__nor2_2 _4128_ (.A(_1705_),
    .B(_1720_),
    .Y(_1724_));
 sky130_fd_sc_hd__o21ai_2 _4129_ (.A1(_1722_),
    .A2(_1724_),
    .B1(_1715_),
    .Y(_1725_));
 sky130_fd_sc_hd__o211ai_2 _4130_ (.A1(_1708_),
    .A2(_1709_),
    .B1(_1723_),
    .C1(_1725_),
    .Y(_1726_));
 sky130_fd_sc_hd__and2b_2 _4131_ (.A_N(out_data_flat[239]),
    .B(out_data_flat[207]),
    .X(_1727_));
 sky130_fd_sc_hd__o22a_2 _4132_ (.A1(_1424_),
    .A2(out_data_flat[207]),
    .B1(out_data_flat[206]),
    .B2(_1425_),
    .X(_1728_));
 sky130_fd_sc_hd__o22a_2 _4133_ (.A1(_1426_),
    .A2(out_data_flat[205]),
    .B1(out_data_flat[204]),
    .B2(_1427_),
    .X(_1729_));
 sky130_fd_sc_hd__a22oi_2 _4134_ (.A1(_1425_),
    .A2(out_data_flat[206]),
    .B1(out_data_flat[205]),
    .B2(_1426_),
    .Y(_1730_));
 sky130_fd_sc_hd__nand2b_2 _4135_ (.A_N(_1729_),
    .B(_1730_),
    .Y(_1731_));
 sky130_fd_sc_hd__a21oi_2 _4136_ (.A1(_1728_),
    .A2(_1731_),
    .B1(_1727_),
    .Y(_1732_));
 sky130_fd_sc_hd__a21oi_2 _4137_ (.A1(_1427_),
    .A2(out_data_flat[204]),
    .B1(_1727_),
    .Y(_1733_));
 sky130_fd_sc_hd__and4_2 _4138_ (.A(_1728_),
    .B(_1729_),
    .C(_1730_),
    .D(_1733_),
    .X(_1734_));
 sky130_fd_sc_hd__nand2b_2 _4139_ (.A_N(out_data_flat[203]),
    .B(out_data_flat[235]),
    .Y(_1735_));
 sky130_fd_sc_hd__nand2b_2 _4140_ (.A_N(out_data_flat[235]),
    .B(out_data_flat[203]),
    .Y(_1736_));
 sky130_fd_sc_hd__nand2b_2 _4141_ (.A_N(out_data_flat[233]),
    .B(out_data_flat[201]),
    .Y(_1737_));
 sky130_fd_sc_hd__xnor2_2 _4142_ (.A(out_data_flat[234]),
    .B(out_data_flat[202]),
    .Y(_1738_));
 sky130_fd_sc_hd__and3_2 _4143_ (.A(_1735_),
    .B(_1736_),
    .C(_1738_),
    .X(_1739_));
 sky130_fd_sc_hd__nand2b_2 _4144_ (.A_N(out_data_flat[201]),
    .B(out_data_flat[233]),
    .Y(_1740_));
 sky130_fd_sc_hd__nand2b_2 _4145_ (.A_N(out_data_flat[200]),
    .B(out_data_flat[232]),
    .Y(_1741_));
 sky130_fd_sc_hd__nand2_2 _4146_ (.A(_1740_),
    .B(_1741_),
    .Y(_1742_));
 sky130_fd_sc_hd__a32o_2 _4147_ (.A1(_1737_),
    .A2(_1739_),
    .A3(_1742_),
    .B1(_1459_),
    .B2(out_data_flat[235]),
    .X(_1743_));
 sky130_fd_sc_hd__a31o_2 _4148_ (.A1(out_data_flat[234]),
    .A2(_1460_),
    .A3(_1736_),
    .B1(_1743_),
    .X(_1744_));
 sky130_fd_sc_hd__and2b_2 _4149_ (.A_N(out_data_flat[193]),
    .B(out_data_flat[225]),
    .X(_1745_));
 sky130_fd_sc_hd__nand2b_2 _4150_ (.A_N(out_data_flat[224]),
    .B(out_data_flat[192]),
    .Y(_1746_));
 sky130_fd_sc_hd__nand2b_2 _4151_ (.A_N(out_data_flat[225]),
    .B(out_data_flat[193]),
    .Y(_1747_));
 sky130_fd_sc_hd__o221a_2 _4152_ (.A1(out_data_flat[226]),
    .A2(_1464_),
    .B1(_1745_),
    .B2(_1746_),
    .C1(_1747_),
    .X(_1748_));
 sky130_fd_sc_hd__a22o_2 _4153_ (.A1(out_data_flat[227]),
    .A2(_1463_),
    .B1(_1464_),
    .B2(out_data_flat[226]),
    .X(_1749_));
 sky130_fd_sc_hd__and2b_2 _4154_ (.A_N(out_data_flat[198]),
    .B(out_data_flat[230]),
    .X(_1750_));
 sky130_fd_sc_hd__nand2b_2 _4155_ (.A_N(out_data_flat[230]),
    .B(out_data_flat[198]),
    .Y(_1751_));
 sky130_fd_sc_hd__nand2b_2 _4156_ (.A_N(out_data_flat[199]),
    .B(out_data_flat[231]),
    .Y(_1752_));
 sky130_fd_sc_hd__nand2b_2 _4157_ (.A_N(out_data_flat[231]),
    .B(out_data_flat[199]),
    .Y(_1753_));
 sky130_fd_sc_hd__and4b_2 _4158_ (.A_N(_1750_),
    .B(_1751_),
    .C(_1752_),
    .D(_1753_),
    .X(_1754_));
 sky130_fd_sc_hd__nand2b_2 _4159_ (.A_N(out_data_flat[197]),
    .B(out_data_flat[229]),
    .Y(_1755_));
 sky130_fd_sc_hd__a21bo_2 _4160_ (.A1(out_data_flat[228]),
    .A2(_1462_),
    .B1_N(_1755_),
    .X(_1756_));
 sky130_fd_sc_hd__nand2b_2 _4161_ (.A_N(out_data_flat[227]),
    .B(out_data_flat[195]),
    .Y(_1757_));
 sky130_fd_sc_hd__nand2b_2 _4162_ (.A_N(out_data_flat[229]),
    .B(out_data_flat[197]),
    .Y(_1758_));
 sky130_fd_sc_hd__xnor2_2 _4163_ (.A(out_data_flat[228]),
    .B(out_data_flat[196]),
    .Y(_1759_));
 sky130_fd_sc_hd__and4_2 _4164_ (.A(_1755_),
    .B(_1757_),
    .C(_1758_),
    .D(_1759_),
    .X(_1760_));
 sky130_fd_sc_hd__o211a_2 _4165_ (.A1(_1748_),
    .A2(_1749_),
    .B1(_1754_),
    .C1(_1760_),
    .X(_1761_));
 sky130_fd_sc_hd__a21bo_2 _4166_ (.A1(_1750_),
    .A2(_1753_),
    .B1_N(_1752_),
    .X(_1762_));
 sky130_fd_sc_hd__a31o_2 _4167_ (.A1(_1754_),
    .A2(_1756_),
    .A3(_1758_),
    .B1(_1762_),
    .X(_1763_));
 sky130_fd_sc_hd__nand2b_2 _4168_ (.A_N(out_data_flat[232]),
    .B(out_data_flat[200]),
    .Y(_1764_));
 sky130_fd_sc_hd__and4_2 _4169_ (.A(_1737_),
    .B(_1740_),
    .C(_1741_),
    .D(_1764_),
    .X(_1765_));
 sky130_fd_sc_hd__o211a_2 _4170_ (.A1(_1761_),
    .A2(_1763_),
    .B1(_1765_),
    .C1(_1734_),
    .X(_1766_));
 sky130_fd_sc_hd__a221o_2 _4171_ (.A1(_1734_),
    .A2(_1744_),
    .B1(_1766_),
    .B2(_1739_),
    .C1(_1732_),
    .X(_1767_));
 sky130_fd_sc_hd__o211a_2 _4172_ (.A1(out_data_flat[240]),
    .A2(_1457_),
    .B1(_1715_),
    .C1(_1721_),
    .X(_1768_));
 sky130_fd_sc_hd__a221o_2 _4173_ (.A1(out_data_flat[255]),
    .A2(_1449_),
    .B1(_1693_),
    .B2(_1694_),
    .C1(\gen_pe[1].pe_inst.sel ),
    .X(_1769_));
 sky130_fd_sc_hd__o32a_2 _4174_ (.A1(_1700_),
    .A2(_1701_),
    .A3(_1703_),
    .B1(_1698_),
    .B2(_1697_),
    .X(_1770_));
 sky130_fd_sc_hd__and2b_2 _4175_ (.A_N(_1770_),
    .B(_1696_),
    .X(_1771_));
 sky130_fd_sc_hd__a211o_2 _4176_ (.A1(_1704_),
    .A2(_1726_),
    .B1(_1769_),
    .C1(_1771_),
    .X(_1772_));
 sky130_fd_sc_hd__and4_2 _4177_ (.A(_1704_),
    .B(_1705_),
    .C(_1767_),
    .D(_1768_),
    .X(_1773_));
 sky130_fd_sc_hd__nor2_2 _4178_ (.A(_1690_),
    .B(_1691_),
    .Y(_1774_));
 sky130_fd_sc_hd__or3_2 _4179_ (.A(_1772_),
    .B(_1773_),
    .C(_1774_),
    .X(_1775_));
 sky130_fd_sc_hd__mux2_1 _4180_ (.A0(out_data_flat[224]),
    .A1(out_data_flat[192]),
    .S(_1775_),
    .X(_0577_));
 sky130_fd_sc_hd__mux2_1 _4181_ (.A0(out_data_flat[225]),
    .A1(out_data_flat[193]),
    .S(_1775_),
    .X(_0588_));
 sky130_fd_sc_hd__mux2_1 _4182_ (.A0(out_data_flat[226]),
    .A1(out_data_flat[194]),
    .S(_1775_),
    .X(_0599_));
 sky130_fd_sc_hd__mux2_1 _4183_ (.A0(out_data_flat[227]),
    .A1(out_data_flat[195]),
    .S(_1775_),
    .X(_0602_));
 sky130_fd_sc_hd__mux2_1 _4184_ (.A0(out_data_flat[228]),
    .A1(out_data_flat[196]),
    .S(_1775_),
    .X(_0603_));
 sky130_fd_sc_hd__mux2_1 _4185_ (.A0(out_data_flat[229]),
    .A1(out_data_flat[197]),
    .S(_1775_),
    .X(_0604_));
 sky130_fd_sc_hd__mux2_1 _4186_ (.A0(out_data_flat[230]),
    .A1(out_data_flat[198]),
    .S(_1775_),
    .X(_0605_));
 sky130_fd_sc_hd__mux2_1 _4187_ (.A0(out_data_flat[231]),
    .A1(out_data_flat[199]),
    .S(_1775_),
    .X(_0606_));
 sky130_fd_sc_hd__mux2_1 _4188_ (.A0(out_data_flat[232]),
    .A1(out_data_flat[200]),
    .S(_1775_),
    .X(_0607_));
 sky130_fd_sc_hd__mux2_1 _4189_ (.A0(out_data_flat[233]),
    .A1(out_data_flat[201]),
    .S(_1775_),
    .X(_0608_));
 sky130_fd_sc_hd__mux2_1 _4190_ (.A0(out_data_flat[234]),
    .A1(out_data_flat[202]),
    .S(_1775_),
    .X(_0578_));
 sky130_fd_sc_hd__mux2_1 _4191_ (.A0(out_data_flat[235]),
    .A1(out_data_flat[203]),
    .S(_1775_),
    .X(_0579_));
 sky130_fd_sc_hd__mux2_1 _4192_ (.A0(out_data_flat[236]),
    .A1(out_data_flat[204]),
    .S(_1775_),
    .X(_0580_));
 sky130_fd_sc_hd__mux2_1 _4193_ (.A0(out_data_flat[237]),
    .A1(out_data_flat[205]),
    .S(_1775_),
    .X(_0581_));
 sky130_fd_sc_hd__mux2_1 _4194_ (.A0(out_data_flat[238]),
    .A1(out_data_flat[206]),
    .S(_1775_),
    .X(_0582_));
 sky130_fd_sc_hd__mux2_1 _4195_ (.A0(out_data_flat[239]),
    .A1(out_data_flat[207]),
    .S(_1775_),
    .X(_0583_));
 sky130_fd_sc_hd__mux2_1 _4196_ (.A0(out_data_flat[240]),
    .A1(out_data_flat[208]),
    .S(_1775_),
    .X(_0584_));
 sky130_fd_sc_hd__mux2_1 _4197_ (.A0(out_data_flat[241]),
    .A1(out_data_flat[209]),
    .S(_1775_),
    .X(_0585_));
 sky130_fd_sc_hd__mux2_1 _4198_ (.A0(out_data_flat[242]),
    .A1(out_data_flat[210]),
    .S(_1775_),
    .X(_0586_));
 sky130_fd_sc_hd__mux2_1 _4199_ (.A0(out_data_flat[243]),
    .A1(out_data_flat[211]),
    .S(_1775_),
    .X(_0587_));
 sky130_fd_sc_hd__mux2_1 _4200_ (.A0(out_data_flat[244]),
    .A1(out_data_flat[212]),
    .S(_1775_),
    .X(_0589_));
 sky130_fd_sc_hd__mux2_1 _4201_ (.A0(out_data_flat[245]),
    .A1(out_data_flat[213]),
    .S(_1775_),
    .X(_0590_));
 sky130_fd_sc_hd__mux2_1 _4202_ (.A0(out_data_flat[246]),
    .A1(out_data_flat[214]),
    .S(_1775_),
    .X(_0591_));
 sky130_fd_sc_hd__mux2_1 _4203_ (.A0(out_data_flat[247]),
    .A1(out_data_flat[215]),
    .S(_1775_),
    .X(_0592_));
 sky130_fd_sc_hd__mux2_1 _4204_ (.A0(out_data_flat[248]),
    .A1(out_data_flat[216]),
    .S(_1775_),
    .X(_0593_));
 sky130_fd_sc_hd__mux2_1 _4205_ (.A0(out_data_flat[249]),
    .A1(out_data_flat[217]),
    .S(_1775_),
    .X(_0594_));
 sky130_fd_sc_hd__mux2_1 _4206_ (.A0(out_data_flat[250]),
    .A1(out_data_flat[218]),
    .S(_1775_),
    .X(_0595_));
 sky130_fd_sc_hd__mux2_1 _4207_ (.A0(out_data_flat[251]),
    .A1(out_data_flat[219]),
    .S(_1775_),
    .X(_0596_));
 sky130_fd_sc_hd__mux2_1 _4208_ (.A0(out_data_flat[252]),
    .A1(out_data_flat[220]),
    .S(_1775_),
    .X(_0597_));
 sky130_fd_sc_hd__mux2_1 _4209_ (.A0(out_data_flat[253]),
    .A1(out_data_flat[221]),
    .S(_1775_),
    .X(_0598_));
 sky130_fd_sc_hd__o21ai_2 _4210_ (.A1(_1772_),
    .A2(_1773_),
    .B1(out_data_flat[222]),
    .Y(_1776_));
 sky130_fd_sc_hd__o21ai_2 _4211_ (.A1(_1418_),
    .A2(_1775_),
    .B1(_1776_),
    .Y(_0600_));
 sky130_fd_sc_hd__o21a_2 _4212_ (.A1(out_data_flat[255]),
    .A2(\gen_pe[1].pe_inst.sel ),
    .B1(out_data_flat[223]),
    .X(_0601_));
 sky130_fd_sc_hd__a22o_2 _4213_ (.A1(_1443_),
    .A2(out_data_flat[77]),
    .B1(out_data_flat[76]),
    .B2(_1444_),
    .X(_1777_));
 sky130_fd_sc_hd__and2b_2 _4214_ (.A_N(out_data_flat[79]),
    .B(out_data_flat[47]),
    .X(_1778_));
 sky130_fd_sc_hd__o21bai_2 _4215_ (.A1(_1444_),
    .A2(out_data_flat[76]),
    .B1_N(_1778_),
    .Y(_1779_));
 sky130_fd_sc_hd__a2bb2o_2 _4216_ (.A1_N(_1475_),
    .A2_N(out_data_flat[46]),
    .B1(_1442_),
    .B2(out_data_flat[79]),
    .X(_1780_));
 sky130_fd_sc_hd__inv_2 _4217_ (.A(_1780_),
    .Y(_1781_));
 sky130_fd_sc_hd__a2bb2o_2 _4218_ (.A1_N(out_data_flat[77]),
    .A2_N(_1443_),
    .B1(out_data_flat[46]),
    .B2(_1475_),
    .X(_1782_));
 sky130_fd_sc_hd__or4_2 _4219_ (.A(_1777_),
    .B(_1779_),
    .C(_1780_),
    .D(_1782_),
    .X(_1783_));
 sky130_fd_sc_hd__o22a_2 _4220_ (.A1(out_data_flat[41]),
    .A2(_1476_),
    .B1(_1477_),
    .B2(out_data_flat[40]),
    .X(_1784_));
 sky130_fd_sc_hd__a22o_2 _4221_ (.A1(_1445_),
    .A2(out_data_flat[75]),
    .B1(out_data_flat[74]),
    .B2(_1446_),
    .X(_1785_));
 sky130_fd_sc_hd__nand2b_2 _4222_ (.A_N(out_data_flat[75]),
    .B(out_data_flat[43]),
    .Y(_1786_));
 sky130_fd_sc_hd__o21ai_2 _4223_ (.A1(_1446_),
    .A2(out_data_flat[74]),
    .B1(_1786_),
    .Y(_1787_));
 sky130_fd_sc_hd__a211o_2 _4224_ (.A1(out_data_flat[41]),
    .A2(_1476_),
    .B1(_1785_),
    .C1(_1787_),
    .X(_1788_));
 sky130_fd_sc_hd__o2bb2a_2 _4225_ (.A1_N(_1785_),
    .A2_N(_1786_),
    .B1(_1788_),
    .B2(_1784_),
    .X(_1789_));
 sky130_fd_sc_hd__o22a_2 _4226_ (.A1(out_data_flat[39]),
    .A2(_1478_),
    .B1(_1479_),
    .B2(out_data_flat[38]),
    .X(_1790_));
 sky130_fd_sc_hd__nor2_2 _4227_ (.A(_1447_),
    .B(out_data_flat[69]),
    .Y(_1791_));
 sky130_fd_sc_hd__o22a_2 _4228_ (.A1(out_data_flat[37]),
    .A2(_1480_),
    .B1(_1481_),
    .B2(out_data_flat[36]),
    .X(_1792_));
 sky130_fd_sc_hd__nand2b_2 _4229_ (.A_N(out_data_flat[33]),
    .B(out_data_flat[65]),
    .Y(_1793_));
 sky130_fd_sc_hd__and2b_2 _4230_ (.A_N(out_data_flat[66]),
    .B(out_data_flat[34]),
    .X(_1794_));
 sky130_fd_sc_hd__and2b_2 _4231_ (.A_N(out_data_flat[65]),
    .B(out_data_flat[33]),
    .X(_1795_));
 sky130_fd_sc_hd__a311o_2 _4232_ (.A1(out_data_flat[32]),
    .A2(_1485_),
    .A3(_1793_),
    .B1(_1794_),
    .C1(_1795_),
    .X(_1796_));
 sky130_fd_sc_hd__o22a_2 _4233_ (.A1(out_data_flat[35]),
    .A2(_1482_),
    .B1(_1483_),
    .B2(out_data_flat[34]),
    .X(_1797_));
 sky130_fd_sc_hd__a22o_2 _4234_ (.A1(out_data_flat[36]),
    .A2(_1481_),
    .B1(_1482_),
    .B2(out_data_flat[35]),
    .X(_1798_));
 sky130_fd_sc_hd__a21o_2 _4235_ (.A1(_1796_),
    .A2(_1797_),
    .B1(_1798_),
    .X(_1799_));
 sky130_fd_sc_hd__a221o_2 _4236_ (.A1(out_data_flat[38]),
    .A2(_1479_),
    .B1(_1792_),
    .B2(_1799_),
    .C1(_1791_),
    .X(_1800_));
 sky130_fd_sc_hd__a221o_2 _4237_ (.A1(out_data_flat[40]),
    .A2(_1477_),
    .B1(_1478_),
    .B2(out_data_flat[39]),
    .C1(_1788_),
    .X(_1801_));
 sky130_fd_sc_hd__nand2b_2 _4238_ (.A_N(_1783_),
    .B(_1784_),
    .Y(_1802_));
 sky130_fd_sc_hd__a211o_2 _4239_ (.A1(_1790_),
    .A2(_1800_),
    .B1(_1801_),
    .C1(_1802_),
    .X(_1803_));
 sky130_fd_sc_hd__or4bb_2 _4240_ (.A(_1782_),
    .B(_1778_),
    .C_N(_1777_),
    .D_N(_1781_),
    .X(_1804_));
 sky130_fd_sc_hd__o221a_2 _4241_ (.A1(_1778_),
    .A2(_1781_),
    .B1(_1783_),
    .B2(_1789_),
    .C1(_1804_),
    .X(_1805_));
 sky130_fd_sc_hd__nor2_2 _4242_ (.A(out_data_flat[63]),
    .B(_1465_),
    .Y(_1806_));
 sky130_fd_sc_hd__nor2_2 _4243_ (.A(_1429_),
    .B(out_data_flat[95]),
    .Y(_1807_));
 sky130_fd_sc_hd__a22o_2 _4244_ (.A1(_1430_),
    .A2(out_data_flat[94]),
    .B1(_1467_),
    .B2(out_data_flat[61]),
    .X(_1808_));
 sky130_fd_sc_hd__a2111o_2 _4245_ (.A1(out_data_flat[62]),
    .A2(_1466_),
    .B1(_1806_),
    .C1(_1807_),
    .D1(_1808_),
    .X(_1809_));
 sky130_fd_sc_hd__xor2_2 _4246_ (.A(out_data_flat[58]),
    .B(out_data_flat[90]),
    .X(_1810_));
 sky130_fd_sc_hd__a221o_2 _4247_ (.A1(out_data_flat[59]),
    .A2(_1469_),
    .B1(_1471_),
    .B2(out_data_flat[57]),
    .C1(_1810_),
    .X(_1811_));
 sky130_fd_sc_hd__o22a_2 _4248_ (.A1(out_data_flat[57]),
    .A2(_1471_),
    .B1(_1472_),
    .B2(out_data_flat[56]),
    .X(_1812_));
 sky130_fd_sc_hd__o221ai_2 _4249_ (.A1(out_data_flat[61]),
    .A2(_1467_),
    .B1(_1468_),
    .B2(out_data_flat[60]),
    .C1(_1812_),
    .Y(_1813_));
 sky130_fd_sc_hd__nor2_2 _4250_ (.A(out_data_flat[59]),
    .B(_1469_),
    .Y(_1814_));
 sky130_fd_sc_hd__a221o_2 _4251_ (.A1(out_data_flat[60]),
    .A2(_1468_),
    .B1(_1472_),
    .B2(out_data_flat[56]),
    .C1(_1814_),
    .X(_1815_));
 sky130_fd_sc_hd__or4_2 _4252_ (.A(_1809_),
    .B(_1811_),
    .C(_1813_),
    .D(_1815_),
    .X(_1816_));
 sky130_fd_sc_hd__xor2_2 _4253_ (.A(out_data_flat[50]),
    .B(out_data_flat[82]),
    .X(_1817_));
 sky130_fd_sc_hd__nor2_2 _4254_ (.A(_1440_),
    .B(out_data_flat[81]),
    .Y(_1818_));
 sky130_fd_sc_hd__nand2b_2 _4255_ (.A_N(out_data_flat[51]),
    .B(out_data_flat[83]),
    .Y(_1819_));
 sky130_fd_sc_hd__and2b_2 _4256_ (.A_N(out_data_flat[83]),
    .B(out_data_flat[51]),
    .X(_1820_));
 sky130_fd_sc_hd__or3b_2 _4257_ (.A(_1820_),
    .B(_1817_),
    .C_N(_1819_),
    .X(_1821_));
 sky130_fd_sc_hd__a22o_2 _4258_ (.A1(_1434_),
    .A2(out_data_flat[87]),
    .B1(out_data_flat[86]),
    .B2(_1435_),
    .X(_1822_));
 sky130_fd_sc_hd__a22o_2 _4259_ (.A1(_1436_),
    .A2(out_data_flat[85]),
    .B1(out_data_flat[84]),
    .B2(_1437_),
    .X(_1823_));
 sky130_fd_sc_hd__and2b_2 _4260_ (.A_N(out_data_flat[87]),
    .B(out_data_flat[55]),
    .X(_1824_));
 sky130_fd_sc_hd__o21bai_2 _4261_ (.A1(_1437_),
    .A2(out_data_flat[84]),
    .B1_N(_1824_),
    .Y(_1825_));
 sky130_fd_sc_hd__o22a_2 _4262_ (.A1(_1435_),
    .A2(out_data_flat[86]),
    .B1(out_data_flat[85]),
    .B2(_1436_),
    .X(_1826_));
 sky130_fd_sc_hd__or4b_2 _4263_ (.A(_1822_),
    .B(_1823_),
    .C(_1825_),
    .D_N(_1826_),
    .X(_1827_));
 sky130_fd_sc_hd__o22a_2 _4264_ (.A1(out_data_flat[49]),
    .A2(_1473_),
    .B1(_1474_),
    .B2(out_data_flat[48]),
    .X(_1828_));
 sky130_fd_sc_hd__nor2_2 _4265_ (.A(_1441_),
    .B(out_data_flat[80]),
    .Y(_1829_));
 sky130_fd_sc_hd__or3b_2 _4266_ (.A(_1827_),
    .B(_1829_),
    .C_N(_1828_),
    .X(_1830_));
 sky130_fd_sc_hd__or4_2 _4267_ (.A(_1816_),
    .B(_1818_),
    .C(_1821_),
    .D(_1830_),
    .X(_1831_));
 sky130_fd_sc_hd__a21o_2 _4268_ (.A1(_1803_),
    .A2(_1805_),
    .B1(_1831_),
    .X(_1832_));
 sky130_fd_sc_hd__or3b_2 _4269_ (.A(out_data_flat[50]),
    .B(_1820_),
    .C_N(out_data_flat[82]),
    .X(_1833_));
 sky130_fd_sc_hd__o311a_2 _4270_ (.A1(_1818_),
    .A2(_1821_),
    .A3(_1828_),
    .B1(_1833_),
    .C1(_1819_),
    .X(_1834_));
 sky130_fd_sc_hd__a21oi_2 _4271_ (.A1(_1823_),
    .A2(_1826_),
    .B1(_1822_),
    .Y(_1835_));
 sky130_fd_sc_hd__o22a_2 _4272_ (.A1(_1827_),
    .A2(_1834_),
    .B1(_1835_),
    .B2(_1824_),
    .X(_1836_));
 sky130_fd_sc_hd__a211o_2 _4273_ (.A1(out_data_flat[59]),
    .A2(_1469_),
    .B1(_1470_),
    .C1(out_data_flat[58]),
    .X(_1837_));
 sky130_fd_sc_hd__o221a_2 _4274_ (.A1(out_data_flat[59]),
    .A2(_1469_),
    .B1(_1811_),
    .B2(_1812_),
    .C1(_1837_),
    .X(_1838_));
 sky130_fd_sc_hd__a21o_2 _4275_ (.A1(out_data_flat[60]),
    .A2(_1468_),
    .B1(_1838_),
    .X(_1839_));
 sky130_fd_sc_hd__o221a_2 _4276_ (.A1(out_data_flat[61]),
    .A2(_1467_),
    .B1(_1468_),
    .B2(out_data_flat[60]),
    .C1(_1839_),
    .X(_1840_));
 sky130_fd_sc_hd__or3b_2 _4277_ (.A(out_data_flat[62]),
    .B(_1807_),
    .C_N(out_data_flat[94]),
    .X(_1841_));
 sky130_fd_sc_hd__o221a_2 _4278_ (.A1(out_data_flat[63]),
    .A2(_1465_),
    .B1(_1816_),
    .B2(_1836_),
    .C1(_1841_),
    .X(_1842_));
 sky130_fd_sc_hd__o211a_2 _4279_ (.A1(_1809_),
    .A2(_1840_),
    .B1(_1842_),
    .C1(\gen_pe[1].pe_inst.sel ),
    .X(_1843_));
 sky130_fd_sc_hd__nand2_2 _4280_ (.A(_1832_),
    .B(_1843_),
    .Y(_1844_));
 sky130_fd_sc_hd__mux2_1 _4281_ (.A0(out_data_flat[32]),
    .A1(out_data_flat[64]),
    .S(_1844_),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _4282_ (.A0(out_data_flat[33]),
    .A1(out_data_flat[65]),
    .S(_1844_),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _4283_ (.A0(out_data_flat[34]),
    .A1(out_data_flat[66]),
    .S(_1844_),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _4284_ (.A0(out_data_flat[35]),
    .A1(out_data_flat[67]),
    .S(_1844_),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _4285_ (.A0(out_data_flat[36]),
    .A1(out_data_flat[68]),
    .S(_1844_),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _4286_ (.A0(out_data_flat[37]),
    .A1(out_data_flat[69]),
    .S(_1844_),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _4287_ (.A0(out_data_flat[38]),
    .A1(out_data_flat[70]),
    .S(_1844_),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _4288_ (.A0(out_data_flat[39]),
    .A1(out_data_flat[71]),
    .S(_1844_),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _4289_ (.A0(out_data_flat[40]),
    .A1(out_data_flat[72]),
    .S(_1844_),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _4290_ (.A0(out_data_flat[41]),
    .A1(out_data_flat[73]),
    .S(_1844_),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _4291_ (.A0(out_data_flat[42]),
    .A1(out_data_flat[74]),
    .S(_1844_),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _4292_ (.A0(out_data_flat[43]),
    .A1(out_data_flat[75]),
    .S(_1844_),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_1 _4293_ (.A0(out_data_flat[44]),
    .A1(out_data_flat[76]),
    .S(_1844_),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _4294_ (.A0(out_data_flat[45]),
    .A1(out_data_flat[77]),
    .S(_1844_),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _4295_ (.A0(out_data_flat[46]),
    .A1(out_data_flat[78]),
    .S(_1844_),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _4296_ (.A0(out_data_flat[47]),
    .A1(out_data_flat[79]),
    .S(_1844_),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _4297_ (.A0(out_data_flat[48]),
    .A1(out_data_flat[80]),
    .S(_1844_),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _4298_ (.A0(out_data_flat[49]),
    .A1(out_data_flat[81]),
    .S(_1844_),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _4299_ (.A0(out_data_flat[50]),
    .A1(out_data_flat[82]),
    .S(_1844_),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _4300_ (.A0(out_data_flat[51]),
    .A1(out_data_flat[83]),
    .S(_1844_),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _4301_ (.A0(out_data_flat[52]),
    .A1(out_data_flat[84]),
    .S(_1844_),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _4302_ (.A0(out_data_flat[53]),
    .A1(out_data_flat[85]),
    .S(_1844_),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _4303_ (.A0(out_data_flat[54]),
    .A1(out_data_flat[86]),
    .S(_1844_),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _4304_ (.A0(out_data_flat[55]),
    .A1(out_data_flat[87]),
    .S(_1844_),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _4305_ (.A0(out_data_flat[56]),
    .A1(out_data_flat[88]),
    .S(_1844_),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _4306_ (.A0(out_data_flat[57]),
    .A1(out_data_flat[89]),
    .S(_1844_),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _4307_ (.A0(out_data_flat[58]),
    .A1(out_data_flat[90]),
    .S(_1844_),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _4308_ (.A0(out_data_flat[59]),
    .A1(out_data_flat[91]),
    .S(_1844_),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _4309_ (.A0(out_data_flat[60]),
    .A1(out_data_flat[92]),
    .S(_1844_),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _4310_ (.A0(out_data_flat[61]),
    .A1(out_data_flat[93]),
    .S(_1844_),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _4311_ (.A0(out_data_flat[62]),
    .A1(out_data_flat[94]),
    .S(_1844_),
    .X(_0312_));
 sky130_fd_sc_hd__a21o_2 _4312_ (.A1(\gen_pe[1].pe_inst.sel ),
    .A2(out_data_flat[63]),
    .B1(out_data_flat[95]),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _4313_ (.A0(out_data_flat[64]),
    .A1(out_data_flat[32]),
    .S(_1844_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _4314_ (.A0(out_data_flat[65]),
    .A1(out_data_flat[33]),
    .S(_1844_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _4315_ (.A0(out_data_flat[66]),
    .A1(out_data_flat[34]),
    .S(_1844_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _4316_ (.A0(out_data_flat[67]),
    .A1(out_data_flat[35]),
    .S(_1844_),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _4317_ (.A0(out_data_flat[68]),
    .A1(out_data_flat[36]),
    .S(_1844_),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _4318_ (.A0(out_data_flat[69]),
    .A1(out_data_flat[37]),
    .S(_1844_),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _4319_ (.A0(out_data_flat[70]),
    .A1(out_data_flat[38]),
    .S(_1844_),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _4320_ (.A0(out_data_flat[71]),
    .A1(out_data_flat[39]),
    .S(_1844_),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _4321_ (.A0(out_data_flat[72]),
    .A1(out_data_flat[40]),
    .S(_1844_),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _4322_ (.A0(out_data_flat[73]),
    .A1(out_data_flat[41]),
    .S(_1844_),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_1 _4323_ (.A0(out_data_flat[74]),
    .A1(out_data_flat[42]),
    .S(_1844_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _4324_ (.A0(out_data_flat[75]),
    .A1(out_data_flat[43]),
    .S(_1844_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _4325_ (.A0(out_data_flat[76]),
    .A1(out_data_flat[44]),
    .S(_1844_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _4326_ (.A0(out_data_flat[77]),
    .A1(out_data_flat[45]),
    .S(_1844_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _4327_ (.A0(out_data_flat[78]),
    .A1(out_data_flat[46]),
    .S(_1844_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _4328_ (.A0(out_data_flat[79]),
    .A1(out_data_flat[47]),
    .S(_1844_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _4329_ (.A0(out_data_flat[80]),
    .A1(out_data_flat[48]),
    .S(_1844_),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _4330_ (.A0(out_data_flat[81]),
    .A1(out_data_flat[49]),
    .S(_1844_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _4331_ (.A0(out_data_flat[82]),
    .A1(out_data_flat[50]),
    .S(_1844_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _4332_ (.A0(out_data_flat[83]),
    .A1(out_data_flat[51]),
    .S(_1844_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _4333_ (.A0(out_data_flat[84]),
    .A1(out_data_flat[52]),
    .S(_1844_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _4334_ (.A0(out_data_flat[85]),
    .A1(out_data_flat[53]),
    .S(_1844_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _4335_ (.A0(out_data_flat[86]),
    .A1(out_data_flat[54]),
    .S(_1844_),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _4336_ (.A0(out_data_flat[87]),
    .A1(out_data_flat[55]),
    .S(_1844_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _4337_ (.A0(out_data_flat[88]),
    .A1(out_data_flat[56]),
    .S(_1844_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _4338_ (.A0(out_data_flat[89]),
    .A1(out_data_flat[57]),
    .S(_1844_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _4339_ (.A0(out_data_flat[90]),
    .A1(out_data_flat[58]),
    .S(_1844_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _4340_ (.A0(out_data_flat[91]),
    .A1(out_data_flat[59]),
    .S(_1844_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _4341_ (.A0(out_data_flat[92]),
    .A1(out_data_flat[60]),
    .S(_1844_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _4342_ (.A0(out_data_flat[93]),
    .A1(out_data_flat[61]),
    .S(_1844_),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _4343_ (.A0(out_data_flat[94]),
    .A1(out_data_flat[62]),
    .S(_1844_),
    .X(_0280_));
 sky130_fd_sc_hd__a21oi_2 _4344_ (.A1(\gen_pe[1].pe_inst.sel ),
    .A2(_1465_),
    .B1(_1429_),
    .Y(_0281_));
 sky130_fd_sc_hd__a22o_2 _4345_ (.A1(out_data_flat[93]),
    .A2(_1488_),
    .B1(_1489_),
    .B2(out_data_flat[92]),
    .X(_1845_));
 sky130_fd_sc_hd__o22a_2 _4346_ (.A1(out_data_flat[94]),
    .A2(_1487_),
    .B1(_1488_),
    .B2(out_data_flat[93]),
    .X(_1846_));
 sky130_fd_sc_hd__o2bb2a_2 _4347_ (.A1_N(_1487_),
    .A2_N(out_data_flat[94]),
    .B1(_1465_),
    .B2(out_data_flat[127]),
    .X(_1847_));
 sky130_fd_sc_hd__and2b_2 _4348_ (.A_N(out_data_flat[95]),
    .B(out_data_flat[127]),
    .X(_1848_));
 sky130_fd_sc_hd__a21oi_2 _4349_ (.A1(_1468_),
    .A2(out_data_flat[124]),
    .B1(_1848_),
    .Y(_1849_));
 sky130_fd_sc_hd__and4b_2 _4350_ (.A_N(_1845_),
    .B(_1846_),
    .C(_1847_),
    .D(_1849_),
    .X(_1850_));
 sky130_fd_sc_hd__nand2_2 _4351_ (.A(out_data_flat[91]),
    .B(_1490_),
    .Y(_1851_));
 sky130_fd_sc_hd__o22a_2 _4352_ (.A1(out_data_flat[91]),
    .A2(_1490_),
    .B1(out_data_flat[122]),
    .B2(_1470_),
    .X(_1852_));
 sky130_fd_sc_hd__o211a_2 _4353_ (.A1(out_data_flat[90]),
    .A2(_1491_),
    .B1(_1851_),
    .C1(_1852_),
    .X(_1853_));
 sky130_fd_sc_hd__o22a_2 _4354_ (.A1(_1471_),
    .A2(out_data_flat[121]),
    .B1(out_data_flat[120]),
    .B2(_1472_),
    .X(_1854_));
 sky130_fd_sc_hd__o21a_2 _4355_ (.A1(out_data_flat[88]),
    .A2(_1493_),
    .B1(_1854_),
    .X(_1855_));
 sky130_fd_sc_hd__o2111a_2 _4356_ (.A1(out_data_flat[89]),
    .A2(_1492_),
    .B1(_1850_),
    .C1(_1853_),
    .D1(_1855_),
    .X(_1856_));
 sky130_fd_sc_hd__and2b_2 _4357_ (.A_N(out_data_flat[118]),
    .B(out_data_flat[86]),
    .X(_1857_));
 sky130_fd_sc_hd__and2b_2 _4358_ (.A_N(out_data_flat[119]),
    .B(out_data_flat[87]),
    .X(_1858_));
 sky130_fd_sc_hd__and2b_2 _4359_ (.A_N(out_data_flat[116]),
    .B(out_data_flat[84]),
    .X(_1859_));
 sky130_fd_sc_hd__a2111o_2 _4360_ (.A1(out_data_flat[85]),
    .A2(_1496_),
    .B1(_1857_),
    .C1(_1858_),
    .D1(_1859_),
    .X(_1860_));
 sky130_fd_sc_hd__nand2b_2 _4361_ (.A_N(out_data_flat[87]),
    .B(out_data_flat[119]),
    .Y(_1861_));
 sky130_fd_sc_hd__o21a_2 _4362_ (.A1(out_data_flat[84]),
    .A2(_1497_),
    .B1(_1861_),
    .X(_1862_));
 sky130_fd_sc_hd__o22a_2 _4363_ (.A1(out_data_flat[86]),
    .A2(_1495_),
    .B1(_1496_),
    .B2(out_data_flat[85]),
    .X(_1863_));
 sky130_fd_sc_hd__and3b_2 _4364_ (.A_N(_1860_),
    .B(_1862_),
    .C(_1863_),
    .X(_1864_));
 sky130_fd_sc_hd__and2b_2 _4365_ (.A_N(out_data_flat[115]),
    .B(out_data_flat[83]),
    .X(_1865_));
 sky130_fd_sc_hd__nand2_2 _4366_ (.A(out_data_flat[82]),
    .B(_1499_),
    .Y(_1866_));
 sky130_fd_sc_hd__o21ba_2 _4367_ (.A1(out_data_flat[82]),
    .A2(_1499_),
    .B1_N(_1865_),
    .X(_1867_));
 sky130_fd_sc_hd__o211a_2 _4368_ (.A1(out_data_flat[83]),
    .A2(_1498_),
    .B1(_1866_),
    .C1(_1867_),
    .X(_1868_));
 sky130_fd_sc_hd__o211a_2 _4369_ (.A1(out_data_flat[81]),
    .A2(_1500_),
    .B1(_1864_),
    .C1(_1868_),
    .X(_1869_));
 sky130_fd_sc_hd__o22a_2 _4370_ (.A1(_1473_),
    .A2(out_data_flat[113]),
    .B1(out_data_flat[112]),
    .B2(_1474_),
    .X(_1870_));
 sky130_fd_sc_hd__inv_2 _4371_ (.A(_1870_),
    .Y(_1871_));
 sky130_fd_sc_hd__o2111a_2 _4372_ (.A1(out_data_flat[80]),
    .A2(_1501_),
    .B1(_1856_),
    .C1(_1869_),
    .D1(_1870_),
    .X(_1872_));
 sky130_fd_sc_hd__and2b_2 _4373_ (.A_N(out_data_flat[111]),
    .B(out_data_flat[79]),
    .X(_1873_));
 sky130_fd_sc_hd__and2b_2 _4374_ (.A_N(out_data_flat[79]),
    .B(out_data_flat[111]),
    .X(_1874_));
 sky130_fd_sc_hd__xor2_2 _4375_ (.A(out_data_flat[78]),
    .B(out_data_flat[110]),
    .X(_1875_));
 sky130_fd_sc_hd__or3_2 _4376_ (.A(_1873_),
    .B(_1874_),
    .C(_1875_),
    .X(_1876_));
 sky130_fd_sc_hd__and2b_2 _4377_ (.A_N(out_data_flat[109]),
    .B(out_data_flat[77]),
    .X(_1877_));
 sky130_fd_sc_hd__and2b_2 _4378_ (.A_N(out_data_flat[108]),
    .B(out_data_flat[76]),
    .X(_1878_));
 sky130_fd_sc_hd__nor2_2 _4379_ (.A(_1877_),
    .B(_1878_),
    .Y(_1879_));
 sky130_fd_sc_hd__and2b_2 _4380_ (.A_N(out_data_flat[77]),
    .B(out_data_flat[109]),
    .X(_1880_));
 sky130_fd_sc_hd__and2b_2 _4381_ (.A_N(out_data_flat[76]),
    .B(out_data_flat[108]),
    .X(_1881_));
 sky130_fd_sc_hd__or4_2 _4382_ (.A(_1877_),
    .B(_1878_),
    .C(_1880_),
    .D(_1881_),
    .X(_1882_));
 sky130_fd_sc_hd__and2b_2 _4383_ (.A_N(out_data_flat[75]),
    .B(out_data_flat[107]),
    .X(_1883_));
 sky130_fd_sc_hd__or3b_2 _4384_ (.A(out_data_flat[106]),
    .B(_1883_),
    .C_N(out_data_flat[74]),
    .X(_1884_));
 sky130_fd_sc_hd__and2b_2 _4385_ (.A_N(out_data_flat[107]),
    .B(out_data_flat[75]),
    .X(_1885_));
 sky130_fd_sc_hd__inv_2 _4386_ (.A(_1885_),
    .Y(_1886_));
 sky130_fd_sc_hd__xor2_2 _4387_ (.A(out_data_flat[74]),
    .B(out_data_flat[106]),
    .X(_1887_));
 sky130_fd_sc_hd__and2b_2 _4388_ (.A_N(out_data_flat[73]),
    .B(out_data_flat[105]),
    .X(_1888_));
 sky130_fd_sc_hd__or4_2 _4389_ (.A(_1883_),
    .B(_1885_),
    .C(_1887_),
    .D(_1888_),
    .X(_1889_));
 sky130_fd_sc_hd__and2b_2 _4390_ (.A_N(out_data_flat[104]),
    .B(out_data_flat[72]),
    .X(_1890_));
 sky130_fd_sc_hd__and2b_2 _4391_ (.A_N(out_data_flat[105]),
    .B(out_data_flat[73]),
    .X(_1891_));
 sky130_fd_sc_hd__and2b_2 _4392_ (.A_N(out_data_flat[72]),
    .B(out_data_flat[104]),
    .X(_1892_));
 sky130_fd_sc_hd__and2b_2 _4393_ (.A_N(out_data_flat[71]),
    .B(out_data_flat[103]),
    .X(_1893_));
 sky130_fd_sc_hd__and2b_2 _4394_ (.A_N(out_data_flat[103]),
    .B(out_data_flat[71]),
    .X(_1894_));
 sky130_fd_sc_hd__o22a_2 _4395_ (.A1(_1480_),
    .A2(out_data_flat[101]),
    .B1(out_data_flat[100]),
    .B2(_1481_),
    .X(_1895_));
 sky130_fd_sc_hd__nor2_2 _4396_ (.A(out_data_flat[69]),
    .B(_1503_),
    .Y(_1896_));
 sky130_fd_sc_hd__or3_2 _4397_ (.A(_1475_),
    .B(out_data_flat[110]),
    .C(_1874_),
    .X(_1897_));
 sky130_fd_sc_hd__and2_2 _4398_ (.A(_1481_),
    .B(out_data_flat[100]),
    .X(_1898_));
 sky130_fd_sc_hd__or3_2 _4399_ (.A(_1890_),
    .B(_1891_),
    .C(_1892_),
    .X(_1899_));
 sky130_fd_sc_hd__or4_2 _4400_ (.A(_1876_),
    .B(_1882_),
    .C(_1889_),
    .D(_1899_),
    .X(_1900_));
 sky130_fd_sc_hd__xor2_2 _4401_ (.A(out_data_flat[70]),
    .B(out_data_flat[102]),
    .X(_1901_));
 sky130_fd_sc_hd__or3_2 _4402_ (.A(_1893_),
    .B(_1894_),
    .C(_1901_),
    .X(_1902_));
 sky130_fd_sc_hd__or4b_2 _4403_ (.A(_1896_),
    .B(_1898_),
    .C(_1902_),
    .D_N(_1895_),
    .X(_1903_));
 sky130_fd_sc_hd__nor2_2 _4404_ (.A(_1900_),
    .B(_1903_),
    .Y(_1904_));
 sky130_fd_sc_hd__nand2b_2 _4405_ (.A_N(out_data_flat[99]),
    .B(out_data_flat[67]),
    .Y(_1905_));
 sky130_fd_sc_hd__nand2b_2 _4406_ (.A_N(out_data_flat[67]),
    .B(out_data_flat[99]),
    .Y(_1906_));
 sky130_fd_sc_hd__xnor2_2 _4407_ (.A(out_data_flat[66]),
    .B(out_data_flat[98]),
    .Y(_1907_));
 sky130_fd_sc_hd__and3_2 _4408_ (.A(_1905_),
    .B(_1906_),
    .C(_1907_),
    .X(_1908_));
 sky130_fd_sc_hd__or2_2 _4409_ (.A(_1484_),
    .B(out_data_flat[97]),
    .X(_1909_));
 sky130_fd_sc_hd__a22o_2 _4410_ (.A1(_1484_),
    .A2(out_data_flat[97]),
    .B1(out_data_flat[96]),
    .B2(_1485_),
    .X(_1910_));
 sky130_fd_sc_hd__a21bo_2 _4411_ (.A1(_1909_),
    .A2(_1910_),
    .B1_N(_1908_),
    .X(_1911_));
 sky130_fd_sc_hd__nand3b_2 _4412_ (.A_N(out_data_flat[98]),
    .B(_1906_),
    .C(out_data_flat[66]),
    .Y(_1912_));
 sky130_fd_sc_hd__a311o_2 _4413_ (.A1(_1905_),
    .A2(_1911_),
    .A3(_1912_),
    .B1(_1903_),
    .C1(_1900_),
    .X(_1913_));
 sky130_fd_sc_hd__o32a_2 _4414_ (.A1(_1895_),
    .A2(_1896_),
    .A3(_1902_),
    .B1(out_data_flat[103]),
    .B2(_1478_),
    .X(_1914_));
 sky130_fd_sc_hd__o31a_2 _4415_ (.A1(_1479_),
    .A2(out_data_flat[102]),
    .A3(_1893_),
    .B1(_1914_),
    .X(_1915_));
 sky130_fd_sc_hd__or3_2 _4416_ (.A(_1876_),
    .B(_1879_),
    .C(_1880_),
    .X(_1916_));
 sky130_fd_sc_hd__o21bai_2 _4417_ (.A1(_1890_),
    .A2(_1891_),
    .B1_N(_1888_),
    .Y(_1917_));
 sky130_fd_sc_hd__o311a_2 _4418_ (.A1(_1883_),
    .A2(_1887_),
    .A3(_1917_),
    .B1(_1884_),
    .C1(_1886_),
    .X(_1918_));
 sky130_fd_sc_hd__o31a_2 _4419_ (.A1(_1876_),
    .A2(_1882_),
    .A3(_1918_),
    .B1(_1916_),
    .X(_1919_));
 sky130_fd_sc_hd__and3b_2 _4420_ (.A_N(_1873_),
    .B(_1897_),
    .C(_1919_),
    .X(_1920_));
 sky130_fd_sc_hd__o21a_2 _4421_ (.A1(_1900_),
    .A2(_1915_),
    .B1(_1913_),
    .X(_1921_));
 sky130_fd_sc_hd__a21bo_2 _4422_ (.A1(_1920_),
    .A2(_1921_),
    .B1_N(_1872_),
    .X(_1922_));
 sky130_fd_sc_hd__o311a_2 _4423_ (.A1(_1857_),
    .A2(_1858_),
    .A3(_1863_),
    .B1(_1861_),
    .C1(_1860_),
    .X(_1923_));
 sky130_fd_sc_hd__o211a_2 _4424_ (.A1(out_data_flat[83]),
    .A2(_1498_),
    .B1(_1499_),
    .C1(out_data_flat[82]),
    .X(_1924_));
 sky130_fd_sc_hd__o21a_2 _4425_ (.A1(_1865_),
    .A2(_1924_),
    .B1(_1864_),
    .X(_1925_));
 sky130_fd_sc_hd__a211o_2 _4426_ (.A1(_1869_),
    .A2(_1871_),
    .B1(_1923_),
    .C1(_1925_),
    .X(_1926_));
 sky130_fd_sc_hd__nand2_2 _4427_ (.A(_1845_),
    .B(_1846_),
    .Y(_1927_));
 sky130_fd_sc_hd__a21o_2 _4428_ (.A1(_1847_),
    .A2(_1927_),
    .B1(_1848_),
    .X(_1928_));
 sky130_fd_sc_hd__o211a_2 _4429_ (.A1(out_data_flat[91]),
    .A2(_1490_),
    .B1(_1491_),
    .C1(out_data_flat[90]),
    .X(_1929_));
 sky130_fd_sc_hd__a21oi_2 _4430_ (.A1(_1471_),
    .A2(out_data_flat[121]),
    .B1(_1854_),
    .Y(_1930_));
 sky130_fd_sc_hd__a221o_2 _4431_ (.A1(out_data_flat[91]),
    .A2(_1490_),
    .B1(_1853_),
    .B2(_1930_),
    .C1(_1929_),
    .X(_1931_));
 sky130_fd_sc_hd__a22oi_2 _4432_ (.A1(_1856_),
    .A2(_1926_),
    .B1(_1931_),
    .B2(_1850_),
    .Y(_1932_));
 sky130_fd_sc_hd__o21a_2 _4433_ (.A1(_1485_),
    .A2(out_data_flat[96]),
    .B1(_1908_),
    .X(_1933_));
 sky130_fd_sc_hd__and3b_2 _4434_ (.A_N(_1910_),
    .B(_1933_),
    .C(_1909_),
    .X(_1934_));
 sky130_fd_sc_hd__a31o_2 _4435_ (.A1(_1872_),
    .A2(_1904_),
    .A3(_1934_),
    .B1(\gen_pe[1].pe_inst.sel ),
    .X(_1935_));
 sky130_fd_sc_hd__a31o_2 _4436_ (.A1(_1922_),
    .A2(_1928_),
    .A3(_1932_),
    .B1(_1935_),
    .X(_1936_));
 sky130_fd_sc_hd__mux2_1 _4437_ (.A0(out_data_flat[96]),
    .A1(out_data_flat[64]),
    .S(_1936_),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _4438_ (.A0(out_data_flat[97]),
    .A1(out_data_flat[65]),
    .S(_1936_),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _4439_ (.A0(out_data_flat[98]),
    .A1(out_data_flat[66]),
    .S(_1936_),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_1 _4440_ (.A0(out_data_flat[99]),
    .A1(out_data_flat[67]),
    .S(_1936_),
    .X(_0346_));
 sky130_fd_sc_hd__mux2_1 _4441_ (.A0(out_data_flat[100]),
    .A1(out_data_flat[68]),
    .S(_1936_),
    .X(_0347_));
 sky130_fd_sc_hd__mux2_1 _4442_ (.A0(out_data_flat[101]),
    .A1(out_data_flat[69]),
    .S(_1936_),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_1 _4443_ (.A0(out_data_flat[102]),
    .A1(out_data_flat[70]),
    .S(_1936_),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_1 _4444_ (.A0(out_data_flat[103]),
    .A1(out_data_flat[71]),
    .S(_1936_),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_1 _4445_ (.A0(out_data_flat[104]),
    .A1(out_data_flat[72]),
    .S(_1936_),
    .X(_0351_));
 sky130_fd_sc_hd__mux2_1 _4446_ (.A0(out_data_flat[105]),
    .A1(out_data_flat[73]),
    .S(_1936_),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_1 _4447_ (.A0(out_data_flat[106]),
    .A1(out_data_flat[74]),
    .S(_1936_),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _4448_ (.A0(out_data_flat[107]),
    .A1(out_data_flat[75]),
    .S(_1936_),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _4449_ (.A0(out_data_flat[108]),
    .A1(out_data_flat[76]),
    .S(_1936_),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_1 _4450_ (.A0(out_data_flat[109]),
    .A1(out_data_flat[77]),
    .S(_1936_),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_1 _4451_ (.A0(out_data_flat[110]),
    .A1(out_data_flat[78]),
    .S(_1936_),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_1 _4452_ (.A0(out_data_flat[111]),
    .A1(out_data_flat[79]),
    .S(_1936_),
    .X(_0327_));
 sky130_fd_sc_hd__mux2_1 _4453_ (.A0(out_data_flat[112]),
    .A1(out_data_flat[80]),
    .S(_1936_),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _4454_ (.A0(out_data_flat[113]),
    .A1(out_data_flat[81]),
    .S(_1936_),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _4455_ (.A0(out_data_flat[114]),
    .A1(out_data_flat[82]),
    .S(_1936_),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _4456_ (.A0(out_data_flat[115]),
    .A1(out_data_flat[83]),
    .S(_1936_),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_1 _4457_ (.A0(out_data_flat[116]),
    .A1(out_data_flat[84]),
    .S(_1936_),
    .X(_0333_));
 sky130_fd_sc_hd__mux2_1 _4458_ (.A0(out_data_flat[117]),
    .A1(out_data_flat[85]),
    .S(_1936_),
    .X(_0334_));
 sky130_fd_sc_hd__mux2_1 _4459_ (.A0(out_data_flat[118]),
    .A1(out_data_flat[86]),
    .S(_1936_),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_1 _4460_ (.A0(out_data_flat[119]),
    .A1(out_data_flat[87]),
    .S(_1936_),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _4461_ (.A0(out_data_flat[120]),
    .A1(out_data_flat[88]),
    .S(_1936_),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _4462_ (.A0(out_data_flat[121]),
    .A1(out_data_flat[89]),
    .S(_1936_),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_1 _4463_ (.A0(out_data_flat[122]),
    .A1(out_data_flat[90]),
    .S(_1936_),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_1 _4464_ (.A0(out_data_flat[123]),
    .A1(out_data_flat[91]),
    .S(_1936_),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _4465_ (.A0(out_data_flat[124]),
    .A1(out_data_flat[92]),
    .S(_1936_),
    .X(_0341_));
 sky130_fd_sc_hd__mux2_1 _4466_ (.A0(out_data_flat[125]),
    .A1(out_data_flat[93]),
    .S(_1936_),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_1 _4467_ (.A0(out_data_flat[126]),
    .A1(out_data_flat[94]),
    .S(_1936_),
    .X(_0344_));
 sky130_fd_sc_hd__o21a_2 _4468_ (.A1(\gen_pe[1].pe_inst.sel ),
    .A2(out_data_flat[127]),
    .B1(out_data_flat[95]),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_1 _4469_ (.A0(out_data_flat[64]),
    .A1(out_data_flat[96]),
    .S(_1936_),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _4470_ (.A0(out_data_flat[65]),
    .A1(out_data_flat[97]),
    .S(_1936_),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_1 _4471_ (.A0(out_data_flat[66]),
    .A1(out_data_flat[98]),
    .S(_1936_),
    .X(_0375_));
 sky130_fd_sc_hd__mux2_1 _4472_ (.A0(out_data_flat[67]),
    .A1(out_data_flat[99]),
    .S(_1936_),
    .X(_0378_));
 sky130_fd_sc_hd__mux2_1 _4473_ (.A0(out_data_flat[68]),
    .A1(out_data_flat[100]),
    .S(_1936_),
    .X(_0379_));
 sky130_fd_sc_hd__mux2_1 _4474_ (.A0(out_data_flat[69]),
    .A1(out_data_flat[101]),
    .S(_1936_),
    .X(_0380_));
 sky130_fd_sc_hd__mux2_1 _4475_ (.A0(out_data_flat[70]),
    .A1(out_data_flat[102]),
    .S(_1936_),
    .X(_0381_));
 sky130_fd_sc_hd__mux2_1 _4476_ (.A0(out_data_flat[71]),
    .A1(out_data_flat[103]),
    .S(_1936_),
    .X(_0382_));
 sky130_fd_sc_hd__mux2_1 _4477_ (.A0(out_data_flat[72]),
    .A1(out_data_flat[104]),
    .S(_1936_),
    .X(_0383_));
 sky130_fd_sc_hd__mux2_1 _4478_ (.A0(out_data_flat[73]),
    .A1(out_data_flat[105]),
    .S(_1936_),
    .X(_0384_));
 sky130_fd_sc_hd__mux2_1 _4479_ (.A0(out_data_flat[74]),
    .A1(out_data_flat[106]),
    .S(_1936_),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _4480_ (.A0(out_data_flat[75]),
    .A1(out_data_flat[107]),
    .S(_1936_),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _4481_ (.A0(out_data_flat[76]),
    .A1(out_data_flat[108]),
    .S(_1936_),
    .X(_0356_));
 sky130_fd_sc_hd__mux2_1 _4482_ (.A0(out_data_flat[77]),
    .A1(out_data_flat[109]),
    .S(_1936_),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_1 _4483_ (.A0(out_data_flat[78]),
    .A1(out_data_flat[110]),
    .S(_1936_),
    .X(_0358_));
 sky130_fd_sc_hd__mux2_1 _4484_ (.A0(out_data_flat[79]),
    .A1(out_data_flat[111]),
    .S(_1936_),
    .X(_0359_));
 sky130_fd_sc_hd__mux2_1 _4485_ (.A0(out_data_flat[80]),
    .A1(out_data_flat[112]),
    .S(_1936_),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_1 _4486_ (.A0(out_data_flat[81]),
    .A1(out_data_flat[113]),
    .S(_1936_),
    .X(_0361_));
 sky130_fd_sc_hd__mux2_1 _4487_ (.A0(out_data_flat[82]),
    .A1(out_data_flat[114]),
    .S(_1936_),
    .X(_0362_));
 sky130_fd_sc_hd__mux2_1 _4488_ (.A0(out_data_flat[83]),
    .A1(out_data_flat[115]),
    .S(_1936_),
    .X(_0363_));
 sky130_fd_sc_hd__mux2_1 _4489_ (.A0(out_data_flat[84]),
    .A1(out_data_flat[116]),
    .S(_1936_),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_1 _4490_ (.A0(out_data_flat[85]),
    .A1(out_data_flat[117]),
    .S(_1936_),
    .X(_0366_));
 sky130_fd_sc_hd__mux2_1 _4491_ (.A0(out_data_flat[86]),
    .A1(out_data_flat[118]),
    .S(_1936_),
    .X(_0367_));
 sky130_fd_sc_hd__mux2_1 _4492_ (.A0(out_data_flat[87]),
    .A1(out_data_flat[119]),
    .S(_1936_),
    .X(_0368_));
 sky130_fd_sc_hd__mux2_1 _4493_ (.A0(out_data_flat[88]),
    .A1(out_data_flat[120]),
    .S(_1936_),
    .X(_0369_));
 sky130_fd_sc_hd__mux2_1 _4494_ (.A0(out_data_flat[89]),
    .A1(out_data_flat[121]),
    .S(_1936_),
    .X(_0370_));
 sky130_fd_sc_hd__mux2_1 _4495_ (.A0(out_data_flat[90]),
    .A1(out_data_flat[122]),
    .S(_1936_),
    .X(_0371_));
 sky130_fd_sc_hd__mux2_1 _4496_ (.A0(out_data_flat[91]),
    .A1(out_data_flat[123]),
    .S(_1936_),
    .X(_0372_));
 sky130_fd_sc_hd__mux2_1 _4497_ (.A0(out_data_flat[92]),
    .A1(out_data_flat[124]),
    .S(_1936_),
    .X(_0373_));
 sky130_fd_sc_hd__mux2_1 _4498_ (.A0(out_data_flat[93]),
    .A1(out_data_flat[125]),
    .S(_1936_),
    .X(_0374_));
 sky130_fd_sc_hd__mux2_1 _4499_ (.A0(out_data_flat[94]),
    .A1(out_data_flat[126]),
    .S(_1936_),
    .X(_0376_));
 sky130_fd_sc_hd__a21o_2 _4500_ (.A1(_1428_),
    .A2(out_data_flat[95]),
    .B1(out_data_flat[127]),
    .X(_0377_));
 sky130_fd_sc_hd__a22o_2 _4501_ (.A1(out_data_flat[217]),
    .A2(_1507_),
    .B1(_1508_),
    .B2(out_data_flat[216]),
    .X(_1937_));
 sky130_fd_sc_hd__o22a_2 _4502_ (.A1(_1449_),
    .A2(out_data_flat[191]),
    .B1(out_data_flat[190]),
    .B2(_1450_),
    .X(_1938_));
 sky130_fd_sc_hd__and2b_2 _4503_ (.A_N(out_data_flat[223]),
    .B(out_data_flat[191]),
    .X(_1939_));
 sky130_fd_sc_hd__a21oi_2 _4504_ (.A1(_1450_),
    .A2(out_data_flat[190]),
    .B1(_1939_),
    .Y(_1940_));
 sky130_fd_sc_hd__o211ai_2 _4505_ (.A1(out_data_flat[221]),
    .A2(_1505_),
    .B1(_1938_),
    .C1(_1940_),
    .Y(_1941_));
 sky130_fd_sc_hd__o22a_2 _4506_ (.A1(_1451_),
    .A2(out_data_flat[189]),
    .B1(out_data_flat[188]),
    .B2(_1452_),
    .X(_1942_));
 sky130_fd_sc_hd__and2b_2 _4507_ (.A_N(out_data_flat[219]),
    .B(out_data_flat[187]),
    .X(_1943_));
 sky130_fd_sc_hd__nor2_2 _4508_ (.A(out_data_flat[220]),
    .B(_1506_),
    .Y(_1944_));
 sky130_fd_sc_hd__and2b_2 _4509_ (.A_N(out_data_flat[187]),
    .B(out_data_flat[219]),
    .X(_1945_));
 sky130_fd_sc_hd__nor2_2 _4510_ (.A(out_data_flat[217]),
    .B(_1507_),
    .Y(_1946_));
 sky130_fd_sc_hd__o221a_2 _4511_ (.A1(_1938_),
    .A2(_1939_),
    .B1(_1941_),
    .B2(_1942_),
    .C1(\gen_pe[1].pe_inst.sel ),
    .X(_1947_));
 sky130_fd_sc_hd__or3b_2 _4512_ (.A(_1941_),
    .B(_1944_),
    .C_N(_1942_),
    .X(_1948_));
 sky130_fd_sc_hd__xor2_2 _4513_ (.A(out_data_flat[218]),
    .B(out_data_flat[186]),
    .X(_1949_));
 sky130_fd_sc_hd__or3_2 _4514_ (.A(_1943_),
    .B(_1945_),
    .C(_1949_),
    .X(_1950_));
 sky130_fd_sc_hd__or3b_2 _4515_ (.A(_1950_),
    .B(_1946_),
    .C_N(_1937_),
    .X(_1951_));
 sky130_fd_sc_hd__or3b_2 _4516_ (.A(out_data_flat[186]),
    .B(_1943_),
    .C_N(out_data_flat[218]),
    .X(_1952_));
 sky130_fd_sc_hd__and3b_2 _4517_ (.A_N(_1945_),
    .B(_1951_),
    .C(_1952_),
    .X(_1953_));
 sky130_fd_sc_hd__o21a_2 _4518_ (.A1(_1948_),
    .A2(_1953_),
    .B1(_1947_),
    .X(_1954_));
 sky130_fd_sc_hd__a2111o_2 _4519_ (.A1(_1453_),
    .A2(out_data_flat[184]),
    .B1(_1937_),
    .C1(_1946_),
    .D1(_1948_),
    .X(_1955_));
 sky130_fd_sc_hd__or2_2 _4520_ (.A(_1950_),
    .B(_1955_),
    .X(_1956_));
 sky130_fd_sc_hd__and2b_2 _4521_ (.A_N(out_data_flat[167]),
    .B(out_data_flat[199]),
    .X(_1957_));
 sky130_fd_sc_hd__and2b_2 _4522_ (.A_N(out_data_flat[166]),
    .B(out_data_flat[198]),
    .X(_1958_));
 sky130_fd_sc_hd__o22a_2 _4523_ (.A1(_1461_),
    .A2(out_data_flat[165]),
    .B1(out_data_flat[164]),
    .B2(_1462_),
    .X(_1959_));
 sky130_fd_sc_hd__nor2_2 _4524_ (.A(out_data_flat[194]),
    .B(_1519_),
    .Y(_1960_));
 sky130_fd_sc_hd__and2b_2 _4525_ (.A_N(out_data_flat[193]),
    .B(out_data_flat[161]),
    .X(_1961_));
 sky130_fd_sc_hd__and2b_2 _4526_ (.A_N(out_data_flat[192]),
    .B(out_data_flat[160]),
    .X(_1962_));
 sky130_fd_sc_hd__nand2b_2 _4527_ (.A_N(out_data_flat[161]),
    .B(out_data_flat[193]),
    .Y(_1963_));
 sky130_fd_sc_hd__o221a_2 _4528_ (.A1(_1464_),
    .A2(out_data_flat[162]),
    .B1(_1961_),
    .B2(_1962_),
    .C1(_1963_),
    .X(_1964_));
 sky130_fd_sc_hd__o22a_2 _4529_ (.A1(_1463_),
    .A2(out_data_flat[163]),
    .B1(_1960_),
    .B2(_1964_),
    .X(_1965_));
 sky130_fd_sc_hd__and2_2 _4530_ (.A(_1463_),
    .B(out_data_flat[163]),
    .X(_1966_));
 sky130_fd_sc_hd__and2b_2 _4531_ (.A_N(out_data_flat[198]),
    .B(out_data_flat[166]),
    .X(_1967_));
 sky130_fd_sc_hd__nand2b_2 _4532_ (.A_N(out_data_flat[206]),
    .B(out_data_flat[174]),
    .Y(_1968_));
 sky130_fd_sc_hd__nor2_2 _4533_ (.A(out_data_flat[205]),
    .B(_1515_),
    .Y(_1969_));
 sky130_fd_sc_hd__nand2b_2 _4534_ (.A_N(out_data_flat[207]),
    .B(out_data_flat[175]),
    .Y(_1970_));
 sky130_fd_sc_hd__and2_2 _4535_ (.A(_1458_),
    .B(out_data_flat[172]),
    .X(_1971_));
 sky130_fd_sc_hd__nand2b_2 _4536_ (.A_N(out_data_flat[175]),
    .B(out_data_flat[207]),
    .Y(_1972_));
 sky130_fd_sc_hd__nand2b_2 _4537_ (.A_N(out_data_flat[174]),
    .B(out_data_flat[206]),
    .Y(_1973_));
 sky130_fd_sc_hd__a2bb2o_2 _4538_ (.A1_N(out_data_flat[172]),
    .A2_N(_1458_),
    .B1(out_data_flat[205]),
    .B2(_1515_),
    .X(_1974_));
 sky130_fd_sc_hd__and4_2 _4539_ (.A(_1968_),
    .B(_1970_),
    .C(_1972_),
    .D(_1973_),
    .X(_1975_));
 sky130_fd_sc_hd__or4b_2 _4540_ (.A(_1969_),
    .B(_1971_),
    .C(_1974_),
    .D_N(_1975_),
    .X(_1976_));
 sky130_fd_sc_hd__nand2b_2 _4541_ (.A_N(out_data_flat[171]),
    .B(out_data_flat[203]),
    .Y(_1977_));
 sky130_fd_sc_hd__and2b_2 _4542_ (.A_N(out_data_flat[203]),
    .B(out_data_flat[171]),
    .X(_1978_));
 sky130_fd_sc_hd__or2_2 _4543_ (.A(out_data_flat[201]),
    .B(_1516_),
    .X(_1979_));
 sky130_fd_sc_hd__xor2_2 _4544_ (.A(out_data_flat[202]),
    .B(out_data_flat[170]),
    .X(_1980_));
 sky130_fd_sc_hd__or3b_2 _4545_ (.A(_1980_),
    .B(_1978_),
    .C_N(_1977_),
    .X(_1981_));
 sky130_fd_sc_hd__a22o_2 _4546_ (.A1(out_data_flat[201]),
    .A2(_1516_),
    .B1(_1517_),
    .B2(out_data_flat[200]),
    .X(_1982_));
 sky130_fd_sc_hd__and2b_2 _4547_ (.A_N(out_data_flat[199]),
    .B(out_data_flat[167]),
    .X(_1983_));
 sky130_fd_sc_hd__nor2_2 _4548_ (.A(out_data_flat[166]),
    .B(_1983_),
    .Y(_1984_));
 sky130_fd_sc_hd__a21oi_2 _4549_ (.A1(out_data_flat[198]),
    .A2(_1984_),
    .B1(_1957_),
    .Y(_1985_));
 sky130_fd_sc_hd__or4_2 _4550_ (.A(_1957_),
    .B(_1958_),
    .C(_1967_),
    .D(_1983_),
    .X(_1986_));
 sky130_fd_sc_hd__a211o_2 _4551_ (.A1(_1461_),
    .A2(out_data_flat[165]),
    .B1(_1959_),
    .C1(_1986_),
    .X(_1987_));
 sky130_fd_sc_hd__a22o_2 _4552_ (.A1(_1461_),
    .A2(out_data_flat[165]),
    .B1(out_data_flat[164]),
    .B2(_1462_),
    .X(_1988_));
 sky130_fd_sc_hd__or4b_2 _4553_ (.A(_1966_),
    .B(_1986_),
    .C(_1988_),
    .D_N(_1959_),
    .X(_1989_));
 sky130_fd_sc_hd__o211a_2 _4554_ (.A1(_1965_),
    .A2(_1989_),
    .B1(_1987_),
    .C1(_1985_),
    .X(_1990_));
 sky130_fd_sc_hd__o21ai_2 _4555_ (.A1(out_data_flat[200]),
    .A2(_1517_),
    .B1(_1979_),
    .Y(_1991_));
 sky130_fd_sc_hd__or4_2 _4556_ (.A(_1976_),
    .B(_1981_),
    .C(_1982_),
    .D(_1991_),
    .X(_1992_));
 sky130_fd_sc_hd__or2_2 _4557_ (.A(_1990_),
    .B(_1992_),
    .X(_1993_));
 sky130_fd_sc_hd__or3_2 _4558_ (.A(_1460_),
    .B(out_data_flat[170]),
    .C(_1978_),
    .X(_1994_));
 sky130_fd_sc_hd__a21bo_2 _4559_ (.A1(_1972_),
    .A2(_1973_),
    .B1_N(_1970_),
    .X(_1995_));
 sky130_fd_sc_hd__nand3b_2 _4560_ (.A_N(_1969_),
    .B(_1974_),
    .C(_1975_),
    .Y(_1996_));
 sky130_fd_sc_hd__nand3b_2 _4561_ (.A_N(_1981_),
    .B(_1982_),
    .C(_1979_),
    .Y(_1997_));
 sky130_fd_sc_hd__a31o_2 _4562_ (.A1(_1977_),
    .A2(_1994_),
    .A3(_1997_),
    .B1(_1976_),
    .X(_1998_));
 sky130_fd_sc_hd__and3_2 _4563_ (.A(_1995_),
    .B(_1996_),
    .C(_1998_),
    .X(_1999_));
 sky130_fd_sc_hd__o2bb2a_2 _4564_ (.A1_N(_1456_),
    .A2_N(out_data_flat[178]),
    .B1(_1513_),
    .B2(out_data_flat[209]),
    .X(_2000_));
 sky130_fd_sc_hd__or2_2 _4565_ (.A(out_data_flat[215]),
    .B(_1509_),
    .X(_2001_));
 sky130_fd_sc_hd__or2_2 _4566_ (.A(out_data_flat[212]),
    .B(_1512_),
    .X(_2002_));
 sky130_fd_sc_hd__nand2_2 _4567_ (.A(_1455_),
    .B(out_data_flat[179]),
    .Y(_2003_));
 sky130_fd_sc_hd__a22oi_2 _4568_ (.A1(out_data_flat[215]),
    .A2(_1509_),
    .B1(_1510_),
    .B2(out_data_flat[214]),
    .Y(_2004_));
 sky130_fd_sc_hd__a22o_2 _4569_ (.A1(out_data_flat[213]),
    .A2(_1511_),
    .B1(_1512_),
    .B2(out_data_flat[212]),
    .X(_2005_));
 sky130_fd_sc_hd__o22a_2 _4570_ (.A1(out_data_flat[214]),
    .A2(_1510_),
    .B1(_1511_),
    .B2(out_data_flat[213]),
    .X(_2006_));
 sky130_fd_sc_hd__and2_2 _4571_ (.A(_2001_),
    .B(_2004_),
    .X(_2007_));
 sky130_fd_sc_hd__and4b_2 _4572_ (.A_N(_2005_),
    .B(_2006_),
    .C(_2007_),
    .D(_2002_),
    .X(_2008_));
 sky130_fd_sc_hd__a22o_2 _4573_ (.A1(out_data_flat[209]),
    .A2(_1513_),
    .B1(_1514_),
    .B2(out_data_flat[208]),
    .X(_2009_));
 sky130_fd_sc_hd__nand2_2 _4574_ (.A(_1457_),
    .B(out_data_flat[176]),
    .Y(_2010_));
 sky130_fd_sc_hd__o22a_2 _4575_ (.A1(_1455_),
    .A2(out_data_flat[179]),
    .B1(out_data_flat[178]),
    .B2(_1456_),
    .X(_2011_));
 sky130_fd_sc_hd__and3b_2 _4576_ (.A_N(_2009_),
    .B(_2010_),
    .C(_2011_),
    .X(_2012_));
 sky130_fd_sc_hd__and4_2 _4577_ (.A(_2000_),
    .B(_2003_),
    .C(_2008_),
    .D(_2012_),
    .X(_2013_));
 sky130_fd_sc_hd__a21bo_2 _4578_ (.A1(_1993_),
    .A2(_1999_),
    .B1_N(_2013_),
    .X(_2014_));
 sky130_fd_sc_hd__a21bo_2 _4579_ (.A1(_2005_),
    .A2(_2006_),
    .B1_N(_2004_),
    .X(_2015_));
 sky130_fd_sc_hd__a21bo_2 _4580_ (.A1(_2000_),
    .A2(_2009_),
    .B1_N(_2011_),
    .X(_2016_));
 sky130_fd_sc_hd__a32o_2 _4581_ (.A1(_2003_),
    .A2(_2008_),
    .A3(_2016_),
    .B1(_2015_),
    .B2(_2001_),
    .X(_2017_));
 sky130_fd_sc_hd__or3b_2 _4582_ (.A(_1950_),
    .B(_1955_),
    .C_N(_2017_),
    .X(_2018_));
 sky130_fd_sc_hd__o211a_2 _4583_ (.A1(_1956_),
    .A2(_2014_),
    .B1(_2018_),
    .C1(_1954_),
    .X(_2019_));
 sky130_fd_sc_hd__mux2_1 _4584_ (.A0(out_data_flat[160]),
    .A1(out_data_flat[192]),
    .S(_2019_),
    .X(_0513_));
 sky130_fd_sc_hd__mux2_1 _4585_ (.A0(out_data_flat[161]),
    .A1(out_data_flat[193]),
    .S(_2019_),
    .X(_0524_));
 sky130_fd_sc_hd__mux2_1 _4586_ (.A0(out_data_flat[162]),
    .A1(out_data_flat[194]),
    .S(_2019_),
    .X(_0535_));
 sky130_fd_sc_hd__mux2_1 _4587_ (.A0(out_data_flat[163]),
    .A1(out_data_flat[195]),
    .S(_2019_),
    .X(_0538_));
 sky130_fd_sc_hd__mux2_1 _4588_ (.A0(out_data_flat[164]),
    .A1(out_data_flat[196]),
    .S(_2019_),
    .X(_0539_));
 sky130_fd_sc_hd__mux2_1 _4589_ (.A0(out_data_flat[165]),
    .A1(out_data_flat[197]),
    .S(_2019_),
    .X(_0540_));
 sky130_fd_sc_hd__mux2_1 _4590_ (.A0(out_data_flat[166]),
    .A1(out_data_flat[198]),
    .S(_2019_),
    .X(_0541_));
 sky130_fd_sc_hd__mux2_1 _4591_ (.A0(out_data_flat[167]),
    .A1(out_data_flat[199]),
    .S(_2019_),
    .X(_0542_));
 sky130_fd_sc_hd__mux2_1 _4592_ (.A0(out_data_flat[168]),
    .A1(out_data_flat[200]),
    .S(_2019_),
    .X(_0543_));
 sky130_fd_sc_hd__mux2_1 _4593_ (.A0(out_data_flat[169]),
    .A1(out_data_flat[201]),
    .S(_2019_),
    .X(_0544_));
 sky130_fd_sc_hd__mux2_1 _4594_ (.A0(out_data_flat[170]),
    .A1(out_data_flat[202]),
    .S(_2019_),
    .X(_0514_));
 sky130_fd_sc_hd__mux2_1 _4595_ (.A0(out_data_flat[171]),
    .A1(out_data_flat[203]),
    .S(_2019_),
    .X(_0515_));
 sky130_fd_sc_hd__mux2_1 _4596_ (.A0(out_data_flat[172]),
    .A1(out_data_flat[204]),
    .S(_2019_),
    .X(_0516_));
 sky130_fd_sc_hd__mux2_1 _4597_ (.A0(out_data_flat[173]),
    .A1(out_data_flat[205]),
    .S(_2019_),
    .X(_0517_));
 sky130_fd_sc_hd__mux2_1 _4598_ (.A0(out_data_flat[174]),
    .A1(out_data_flat[206]),
    .S(_2019_),
    .X(_0518_));
 sky130_fd_sc_hd__mux2_1 _4599_ (.A0(out_data_flat[175]),
    .A1(out_data_flat[207]),
    .S(_2019_),
    .X(_0519_));
 sky130_fd_sc_hd__mux2_1 _4600_ (.A0(out_data_flat[176]),
    .A1(out_data_flat[208]),
    .S(_2019_),
    .X(_0520_));
 sky130_fd_sc_hd__mux2_1 _4601_ (.A0(out_data_flat[177]),
    .A1(out_data_flat[209]),
    .S(_2019_),
    .X(_0521_));
 sky130_fd_sc_hd__mux2_1 _4602_ (.A0(out_data_flat[178]),
    .A1(out_data_flat[210]),
    .S(_2019_),
    .X(_0522_));
 sky130_fd_sc_hd__mux2_1 _4603_ (.A0(out_data_flat[179]),
    .A1(out_data_flat[211]),
    .S(_2019_),
    .X(_0523_));
 sky130_fd_sc_hd__mux2_1 _4604_ (.A0(out_data_flat[180]),
    .A1(out_data_flat[212]),
    .S(_2019_),
    .X(_0525_));
 sky130_fd_sc_hd__mux2_1 _4605_ (.A0(out_data_flat[181]),
    .A1(out_data_flat[213]),
    .S(_2019_),
    .X(_0526_));
 sky130_fd_sc_hd__mux2_1 _4606_ (.A0(out_data_flat[182]),
    .A1(out_data_flat[214]),
    .S(_2019_),
    .X(_0527_));
 sky130_fd_sc_hd__mux2_1 _4607_ (.A0(out_data_flat[183]),
    .A1(out_data_flat[215]),
    .S(_2019_),
    .X(_0528_));
 sky130_fd_sc_hd__mux2_1 _4608_ (.A0(out_data_flat[184]),
    .A1(out_data_flat[216]),
    .S(_2019_),
    .X(_0529_));
 sky130_fd_sc_hd__mux2_1 _4609_ (.A0(out_data_flat[185]),
    .A1(out_data_flat[217]),
    .S(_2019_),
    .X(_0530_));
 sky130_fd_sc_hd__mux2_1 _4610_ (.A0(out_data_flat[186]),
    .A1(out_data_flat[218]),
    .S(_2019_),
    .X(_0531_));
 sky130_fd_sc_hd__mux2_1 _4611_ (.A0(out_data_flat[187]),
    .A1(out_data_flat[219]),
    .S(_2019_),
    .X(_0532_));
 sky130_fd_sc_hd__mux2_1 _4612_ (.A0(out_data_flat[188]),
    .A1(out_data_flat[220]),
    .S(_2019_),
    .X(_0533_));
 sky130_fd_sc_hd__mux2_1 _4613_ (.A0(out_data_flat[189]),
    .A1(out_data_flat[221]),
    .S(_2019_),
    .X(_0534_));
 sky130_fd_sc_hd__mux2_1 _4614_ (.A0(out_data_flat[190]),
    .A1(out_data_flat[222]),
    .S(_2019_),
    .X(_0536_));
 sky130_fd_sc_hd__o21a_2 _4615_ (.A1(_1428_),
    .A2(out_data_flat[223]),
    .B1(out_data_flat[191]),
    .X(_0537_));
 sky130_fd_sc_hd__mux2_1 _4616_ (.A0(out_data_flat[192]),
    .A1(out_data_flat[160]),
    .S(_2019_),
    .X(_0545_));
 sky130_fd_sc_hd__mux2_1 _4617_ (.A0(out_data_flat[193]),
    .A1(out_data_flat[161]),
    .S(_2019_),
    .X(_0556_));
 sky130_fd_sc_hd__mux2_1 _4618_ (.A0(out_data_flat[194]),
    .A1(out_data_flat[162]),
    .S(_2019_),
    .X(_0567_));
 sky130_fd_sc_hd__mux2_1 _4619_ (.A0(out_data_flat[195]),
    .A1(out_data_flat[163]),
    .S(_2019_),
    .X(_0570_));
 sky130_fd_sc_hd__mux2_1 _4620_ (.A0(out_data_flat[196]),
    .A1(out_data_flat[164]),
    .S(_2019_),
    .X(_0571_));
 sky130_fd_sc_hd__mux2_1 _4621_ (.A0(out_data_flat[197]),
    .A1(out_data_flat[165]),
    .S(_2019_),
    .X(_0572_));
 sky130_fd_sc_hd__mux2_1 _4622_ (.A0(out_data_flat[198]),
    .A1(out_data_flat[166]),
    .S(_2019_),
    .X(_0573_));
 sky130_fd_sc_hd__mux2_1 _4623_ (.A0(out_data_flat[199]),
    .A1(out_data_flat[167]),
    .S(_2019_),
    .X(_0574_));
 sky130_fd_sc_hd__mux2_1 _4624_ (.A0(out_data_flat[200]),
    .A1(out_data_flat[168]),
    .S(_2019_),
    .X(_0575_));
 sky130_fd_sc_hd__mux2_1 _4625_ (.A0(out_data_flat[201]),
    .A1(out_data_flat[169]),
    .S(_2019_),
    .X(_0576_));
 sky130_fd_sc_hd__mux2_1 _4626_ (.A0(out_data_flat[202]),
    .A1(out_data_flat[170]),
    .S(_2019_),
    .X(_0546_));
 sky130_fd_sc_hd__mux2_1 _4627_ (.A0(out_data_flat[203]),
    .A1(out_data_flat[171]),
    .S(_2019_),
    .X(_0547_));
 sky130_fd_sc_hd__mux2_1 _4628_ (.A0(out_data_flat[204]),
    .A1(out_data_flat[172]),
    .S(_2019_),
    .X(_0548_));
 sky130_fd_sc_hd__mux2_1 _4629_ (.A0(out_data_flat[205]),
    .A1(out_data_flat[173]),
    .S(_2019_),
    .X(_0549_));
 sky130_fd_sc_hd__mux2_1 _4630_ (.A0(out_data_flat[206]),
    .A1(out_data_flat[174]),
    .S(_2019_),
    .X(_0550_));
 sky130_fd_sc_hd__mux2_1 _4631_ (.A0(out_data_flat[207]),
    .A1(out_data_flat[175]),
    .S(_2019_),
    .X(_0551_));
 sky130_fd_sc_hd__mux2_1 _4632_ (.A0(out_data_flat[208]),
    .A1(out_data_flat[176]),
    .S(_2019_),
    .X(_0552_));
 sky130_fd_sc_hd__mux2_1 _4633_ (.A0(out_data_flat[209]),
    .A1(out_data_flat[177]),
    .S(_2019_),
    .X(_0553_));
 sky130_fd_sc_hd__mux2_1 _4634_ (.A0(out_data_flat[210]),
    .A1(out_data_flat[178]),
    .S(_2019_),
    .X(_0554_));
 sky130_fd_sc_hd__mux2_1 _4635_ (.A0(out_data_flat[211]),
    .A1(out_data_flat[179]),
    .S(_2019_),
    .X(_0555_));
 sky130_fd_sc_hd__mux2_1 _4636_ (.A0(out_data_flat[212]),
    .A1(out_data_flat[180]),
    .S(_2019_),
    .X(_0557_));
 sky130_fd_sc_hd__mux2_1 _4637_ (.A0(out_data_flat[213]),
    .A1(out_data_flat[181]),
    .S(_2019_),
    .X(_0558_));
 sky130_fd_sc_hd__mux2_1 _4638_ (.A0(out_data_flat[214]),
    .A1(out_data_flat[182]),
    .S(_2019_),
    .X(_0559_));
 sky130_fd_sc_hd__mux2_1 _4639_ (.A0(out_data_flat[215]),
    .A1(out_data_flat[183]),
    .S(_2019_),
    .X(_0560_));
 sky130_fd_sc_hd__mux2_1 _4640_ (.A0(out_data_flat[216]),
    .A1(out_data_flat[184]),
    .S(_2019_),
    .X(_0561_));
 sky130_fd_sc_hd__mux2_1 _4641_ (.A0(out_data_flat[217]),
    .A1(out_data_flat[185]),
    .S(_2019_),
    .X(_0562_));
 sky130_fd_sc_hd__mux2_1 _4642_ (.A0(out_data_flat[218]),
    .A1(out_data_flat[186]),
    .S(_2019_),
    .X(_0563_));
 sky130_fd_sc_hd__mux2_1 _4643_ (.A0(out_data_flat[219]),
    .A1(out_data_flat[187]),
    .S(_2019_),
    .X(_0564_));
 sky130_fd_sc_hd__mux2_1 _4644_ (.A0(out_data_flat[220]),
    .A1(out_data_flat[188]),
    .S(_2019_),
    .X(_0565_));
 sky130_fd_sc_hd__mux2_1 _4645_ (.A0(out_data_flat[221]),
    .A1(out_data_flat[189]),
    .S(_2019_),
    .X(_0566_));
 sky130_fd_sc_hd__mux2_1 _4646_ (.A0(out_data_flat[222]),
    .A1(out_data_flat[190]),
    .S(_2019_),
    .X(_0568_));
 sky130_fd_sc_hd__a21o_2 _4647_ (.A1(\gen_pe[1].pe_inst.sel ),
    .A2(out_data_flat[191]),
    .B1(out_data_flat[223]),
    .X(_0569_));
 sky130_fd_sc_hd__and2_2 _4648_ (.A(out_data_flat[187]),
    .B(_1523_),
    .X(_2020_));
 sky130_fd_sc_hd__nor2_2 _4649_ (.A(_1507_),
    .B(out_data_flat[153]),
    .Y(_2021_));
 sky130_fd_sc_hd__or2_2 _4650_ (.A(out_data_flat[187]),
    .B(_1523_),
    .X(_2022_));
 sky130_fd_sc_hd__xor2_2 _4651_ (.A(out_data_flat[186]),
    .B(out_data_flat[154]),
    .X(_2023_));
 sky130_fd_sc_hd__or4b_2 _4652_ (.A(_2020_),
    .B(_2021_),
    .C(_2023_),
    .D_N(_2022_),
    .X(_2024_));
 sky130_fd_sc_hd__a2bb2o_2 _4653_ (.A1_N(out_data_flat[191]),
    .A2_N(_1521_),
    .B1(out_data_flat[158]),
    .B2(_1504_),
    .X(_2025_));
 sky130_fd_sc_hd__a22o_2 _4654_ (.A1(_1505_),
    .A2(out_data_flat[157]),
    .B1(out_data_flat[156]),
    .B2(_1506_),
    .X(_2026_));
 sky130_fd_sc_hd__and2b_2 _4655_ (.A_N(out_data_flat[159]),
    .B(out_data_flat[191]),
    .X(_2027_));
 sky130_fd_sc_hd__a21o_2 _4656_ (.A1(out_data_flat[188]),
    .A2(_1522_),
    .B1(_2027_),
    .X(_2028_));
 sky130_fd_sc_hd__o22a_2 _4657_ (.A1(_1504_),
    .A2(out_data_flat[158]),
    .B1(out_data_flat[157]),
    .B2(_1505_),
    .X(_2029_));
 sky130_fd_sc_hd__or4b_2 _4658_ (.A(_2025_),
    .B(_2026_),
    .C(_2028_),
    .D_N(_2029_),
    .X(_2030_));
 sky130_fd_sc_hd__a22o_2 _4659_ (.A1(_1507_),
    .A2(out_data_flat[153]),
    .B1(out_data_flat[152]),
    .B2(_1508_),
    .X(_2031_));
 sky130_fd_sc_hd__a2111o_2 _4660_ (.A1(out_data_flat[184]),
    .A2(_1524_),
    .B1(_2024_),
    .C1(_2030_),
    .D1(_2031_),
    .X(_2032_));
 sky130_fd_sc_hd__o22a_2 _4661_ (.A1(out_data_flat[177]),
    .A2(_1527_),
    .B1(_1528_),
    .B2(out_data_flat[176]),
    .X(_2033_));
 sky130_fd_sc_hd__o21ai_2 _4662_ (.A1(_1514_),
    .A2(out_data_flat[144]),
    .B1(_2033_),
    .Y(_2034_));
 sky130_fd_sc_hd__nand2b_2 _4663_ (.A_N(out_data_flat[183]),
    .B(out_data_flat[151]),
    .Y(_2035_));
 sky130_fd_sc_hd__nand2b_2 _4664_ (.A_N(out_data_flat[182]),
    .B(out_data_flat[150]),
    .Y(_2036_));
 sky130_fd_sc_hd__nand2b_2 _4665_ (.A_N(out_data_flat[181]),
    .B(out_data_flat[149]),
    .Y(_2037_));
 sky130_fd_sc_hd__o2111a_2 _4666_ (.A1(out_data_flat[180]),
    .A2(_1526_),
    .B1(_2035_),
    .C1(_2036_),
    .D1(_2037_),
    .X(_2038_));
 sky130_fd_sc_hd__nor2_2 _4667_ (.A(_1512_),
    .B(out_data_flat[148]),
    .Y(_2039_));
 sky130_fd_sc_hd__nor2_2 _4668_ (.A(_1509_),
    .B(out_data_flat[151]),
    .Y(_2040_));
 sky130_fd_sc_hd__o22ai_2 _4669_ (.A1(_1510_),
    .A2(out_data_flat[150]),
    .B1(out_data_flat[149]),
    .B2(_1511_),
    .Y(_2041_));
 sky130_fd_sc_hd__or4b_2 _4670_ (.A(_2039_),
    .B(_2040_),
    .C(_2041_),
    .D_N(_2038_),
    .X(_2042_));
 sky130_fd_sc_hd__and2b_2 _4671_ (.A_N(out_data_flat[147]),
    .B(out_data_flat[179]),
    .X(_2043_));
 sky130_fd_sc_hd__nand2b_2 _4672_ (.A_N(out_data_flat[179]),
    .B(out_data_flat[147]),
    .Y(_2044_));
 sky130_fd_sc_hd__nor2_2 _4673_ (.A(_1513_),
    .B(out_data_flat[145]),
    .Y(_2045_));
 sky130_fd_sc_hd__xor2_2 _4674_ (.A(out_data_flat[178]),
    .B(out_data_flat[146]),
    .X(_2046_));
 sky130_fd_sc_hd__or3b_2 _4675_ (.A(_2043_),
    .B(_2046_),
    .C_N(_2044_),
    .X(_2047_));
 sky130_fd_sc_hd__or4_2 _4676_ (.A(_2034_),
    .B(_2042_),
    .C(_2045_),
    .D(_2047_),
    .X(_2048_));
 sky130_fd_sc_hd__or2_2 _4677_ (.A(_2032_),
    .B(_2048_),
    .X(_2049_));
 sky130_fd_sc_hd__and2b_2 _4678_ (.A_N(out_data_flat[175]),
    .B(out_data_flat[143]),
    .X(_2050_));
 sky130_fd_sc_hd__and2b_2 _4679_ (.A_N(out_data_flat[174]),
    .B(out_data_flat[142]),
    .X(_2051_));
 sky130_fd_sc_hd__nor2_2 _4680_ (.A(_2050_),
    .B(_2051_),
    .Y(_2052_));
 sky130_fd_sc_hd__a22o_2 _4681_ (.A1(out_data_flat[174]),
    .A2(_1529_),
    .B1(_1530_),
    .B2(out_data_flat[173]),
    .X(_2053_));
 sky130_fd_sc_hd__and2b_2 _4682_ (.A_N(out_data_flat[172]),
    .B(out_data_flat[140]),
    .X(_2054_));
 sky130_fd_sc_hd__a2111o_2 _4683_ (.A1(_1515_),
    .A2(out_data_flat[141]),
    .B1(_2050_),
    .C1(_2051_),
    .D1(_2054_),
    .X(_2055_));
 sky130_fd_sc_hd__and2b_2 _4684_ (.A_N(out_data_flat[143]),
    .B(out_data_flat[175]),
    .X(_2056_));
 sky130_fd_sc_hd__a21oi_2 _4685_ (.A1(_2052_),
    .A2(_2053_),
    .B1(_2056_),
    .Y(_2057_));
 sky130_fd_sc_hd__a21o_2 _4686_ (.A1(out_data_flat[172]),
    .A2(_1531_),
    .B1(_2056_),
    .X(_2058_));
 sky130_fd_sc_hd__or3_2 _4687_ (.A(_2053_),
    .B(_2055_),
    .C(_2058_),
    .X(_2059_));
 sky130_fd_sc_hd__and2b_2 _4688_ (.A_N(out_data_flat[139]),
    .B(out_data_flat[171]),
    .X(_2060_));
 sky130_fd_sc_hd__and2b_2 _4689_ (.A_N(out_data_flat[171]),
    .B(out_data_flat[139]),
    .X(_2061_));
 sky130_fd_sc_hd__or3_2 _4690_ (.A(out_data_flat[170]),
    .B(_1533_),
    .C(_2060_),
    .X(_2062_));
 sky130_fd_sc_hd__and2b_2 _4691_ (.A_N(_2061_),
    .B(_2062_),
    .X(_2063_));
 sky130_fd_sc_hd__o2bb2a_2 _4692_ (.A1_N(_2055_),
    .A2_N(_2057_),
    .B1(_2059_),
    .B2(_2063_),
    .X(_2064_));
 sky130_fd_sc_hd__xor2_2 _4693_ (.A(out_data_flat[170]),
    .B(out_data_flat[138]),
    .X(_2065_));
 sky130_fd_sc_hd__a2111o_2 _4694_ (.A1(out_data_flat[169]),
    .A2(_1534_),
    .B1(_2060_),
    .C1(_2061_),
    .D1(_2065_),
    .X(_2066_));
 sky130_fd_sc_hd__or4_2 _4695_ (.A(_2053_),
    .B(_2055_),
    .C(_2058_),
    .D(_2066_),
    .X(_2067_));
 sky130_fd_sc_hd__o22a_2 _4696_ (.A1(out_data_flat[169]),
    .A2(_1534_),
    .B1(_1535_),
    .B2(out_data_flat[168]),
    .X(_2068_));
 sky130_fd_sc_hd__and2_2 _4697_ (.A(out_data_flat[167]),
    .B(_1536_),
    .X(_2069_));
 sky130_fd_sc_hd__o22ai_2 _4698_ (.A1(out_data_flat[167]),
    .A2(_1536_),
    .B1(_1537_),
    .B2(out_data_flat[166]),
    .Y(_2070_));
 sky130_fd_sc_hd__a2bb2o_2 _4699_ (.A1_N(_1538_),
    .A2_N(out_data_flat[164]),
    .B1(_1518_),
    .B2(out_data_flat[133]),
    .X(_2071_));
 sky130_fd_sc_hd__and2b_2 _4700_ (.A_N(out_data_flat[134]),
    .B(out_data_flat[166]),
    .X(_2072_));
 sky130_fd_sc_hd__and2b_2 _4701_ (.A_N(out_data_flat[133]),
    .B(out_data_flat[165]),
    .X(_2073_));
 sky130_fd_sc_hd__nor2_2 _4702_ (.A(_2072_),
    .B(_2073_),
    .Y(_2074_));
 sky130_fd_sc_hd__a21oi_2 _4703_ (.A1(_2071_),
    .A2(_2074_),
    .B1(_2070_),
    .Y(_2075_));
 sky130_fd_sc_hd__or3_2 _4704_ (.A(_2069_),
    .B(_2070_),
    .C(_2072_),
    .X(_2076_));
 sky130_fd_sc_hd__or2_2 _4705_ (.A(_2069_),
    .B(_2075_),
    .X(_2077_));
 sky130_fd_sc_hd__and2_2 _4706_ (.A(out_data_flat[163]),
    .B(_1539_),
    .X(_2078_));
 sky130_fd_sc_hd__a2bb2o_2 _4707_ (.A1_N(out_data_flat[163]),
    .A2_N(_1539_),
    .B1(_1540_),
    .B2(out_data_flat[162]),
    .X(_2079_));
 sky130_fd_sc_hd__a211o_2 _4708_ (.A1(_1519_),
    .A2(out_data_flat[130]),
    .B1(_2078_),
    .C1(_2079_),
    .X(_2080_));
 sky130_fd_sc_hd__xor2_2 _4709_ (.A(out_data_flat[161]),
    .B(out_data_flat[129]),
    .X(_2081_));
 sky130_fd_sc_hd__a21o_2 _4710_ (.A1(out_data_flat[160]),
    .A2(_1542_),
    .B1(_2081_),
    .X(_2082_));
 sky130_fd_sc_hd__o21a_2 _4711_ (.A1(out_data_flat[161]),
    .A2(_1541_),
    .B1(_2082_),
    .X(_2083_));
 sky130_fd_sc_hd__or3_2 _4712_ (.A(out_data_flat[162]),
    .B(_1540_),
    .C(_2078_),
    .X(_2084_));
 sky130_fd_sc_hd__o221a_2 _4713_ (.A1(out_data_flat[163]),
    .A2(_1539_),
    .B1(_2080_),
    .B2(_2083_),
    .C1(_2084_),
    .X(_2085_));
 sky130_fd_sc_hd__nand2_2 _4714_ (.A(out_data_flat[164]),
    .B(_1538_),
    .Y(_2086_));
 sky130_fd_sc_hd__or3_2 _4715_ (.A(_2071_),
    .B(_2073_),
    .C(_2076_),
    .X(_2087_));
 sky130_fd_sc_hd__o21ai_2 _4716_ (.A1(_1517_),
    .A2(out_data_flat[136]),
    .B1(_2068_),
    .Y(_2088_));
 sky130_fd_sc_hd__or2_2 _4717_ (.A(_2067_),
    .B(_2088_),
    .X(_2089_));
 sky130_fd_sc_hd__or4b_2 _4718_ (.A(_2073_),
    .B(_2076_),
    .C(_2089_),
    .D_N(_2086_),
    .X(_2090_));
 sky130_fd_sc_hd__or4b_2 _4719_ (.A(_2085_),
    .B(_2087_),
    .C(_2089_),
    .D_N(_2086_),
    .X(_2091_));
 sky130_fd_sc_hd__o221a_2 _4720_ (.A1(_2067_),
    .A2(_2068_),
    .B1(_2077_),
    .B2(_2089_),
    .C1(_2064_),
    .X(_2092_));
 sky130_fd_sc_hd__a21o_2 _4721_ (.A1(_2091_),
    .A2(_2092_),
    .B1(_2049_),
    .X(_2093_));
 sky130_fd_sc_hd__a311o_2 _4722_ (.A1(_2035_),
    .A2(_2036_),
    .A3(_2041_),
    .B1(_2040_),
    .C1(_2038_),
    .X(_2094_));
 sky130_fd_sc_hd__or3b_2 _4723_ (.A(out_data_flat[178]),
    .B(_2043_),
    .C_N(out_data_flat[146]),
    .X(_2095_));
 sky130_fd_sc_hd__or3_2 _4724_ (.A(_2033_),
    .B(_2045_),
    .C(_2047_),
    .X(_2096_));
 sky130_fd_sc_hd__a31o_2 _4725_ (.A1(_2044_),
    .A2(_2095_),
    .A3(_2096_),
    .B1(_2042_),
    .X(_2097_));
 sky130_fd_sc_hd__a21o_2 _4726_ (.A1(_2094_),
    .A2(_2097_),
    .B1(_2032_),
    .X(_2098_));
 sky130_fd_sc_hd__nand2b_2 _4727_ (.A_N(_2024_),
    .B(_2031_),
    .Y(_2099_));
 sky130_fd_sc_hd__or3b_2 _4728_ (.A(out_data_flat[186]),
    .B(_2020_),
    .C_N(out_data_flat[154]),
    .X(_2100_));
 sky130_fd_sc_hd__a31o_2 _4729_ (.A1(_2022_),
    .A2(_2099_),
    .A3(_2100_),
    .B1(_2030_),
    .X(_2101_));
 sky130_fd_sc_hd__a21oi_2 _4730_ (.A1(_2026_),
    .A2(_2029_),
    .B1(_2025_),
    .Y(_2102_));
 sky130_fd_sc_hd__o211a_2 _4731_ (.A1(_2027_),
    .A2(_2102_),
    .B1(_2101_),
    .C1(_2098_),
    .X(_2103_));
 sky130_fd_sc_hd__a211o_2 _4732_ (.A1(_1520_),
    .A2(out_data_flat[128]),
    .B1(_2080_),
    .C1(_2082_),
    .X(_2104_));
 sky130_fd_sc_hd__nor4_2 _4733_ (.A(_2049_),
    .B(_2071_),
    .C(_2090_),
    .D(_2104_),
    .Y(_2105_));
 sky130_fd_sc_hd__a211o_2 _4734_ (.A1(_2093_),
    .A2(_2103_),
    .B1(_2105_),
    .C1(\gen_pe[1].pe_inst.sel ),
    .X(_2106_));
 sky130_fd_sc_hd__mux2_1 _4735_ (.A0(out_data_flat[160]),
    .A1(out_data_flat[128]),
    .S(_2106_),
    .X(_0449_));
 sky130_fd_sc_hd__mux2_1 _4736_ (.A0(out_data_flat[161]),
    .A1(out_data_flat[129]),
    .S(_2106_),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_1 _4737_ (.A0(out_data_flat[162]),
    .A1(out_data_flat[130]),
    .S(_2106_),
    .X(_0471_));
 sky130_fd_sc_hd__mux2_1 _4738_ (.A0(out_data_flat[163]),
    .A1(out_data_flat[131]),
    .S(_2106_),
    .X(_0474_));
 sky130_fd_sc_hd__mux2_1 _4739_ (.A0(out_data_flat[164]),
    .A1(out_data_flat[132]),
    .S(_2106_),
    .X(_0475_));
 sky130_fd_sc_hd__mux2_1 _4740_ (.A0(out_data_flat[165]),
    .A1(out_data_flat[133]),
    .S(_2106_),
    .X(_0476_));
 sky130_fd_sc_hd__mux2_1 _4741_ (.A0(out_data_flat[166]),
    .A1(out_data_flat[134]),
    .S(_2106_),
    .X(_0477_));
 sky130_fd_sc_hd__dfrtp_2 _4742_ (.CLK(clk),
    .D(_0115_),
    .RESET_B(_0641_),
    .Q(out_data_flat[155]));
 sky130_fd_sc_hd__dfrtp_2 _4743_ (.CLK(clk),
    .D(_0116_),
    .RESET_B(_0642_),
    .Q(out_data_flat[156]));
 sky130_fd_sc_hd__dfrtp_2 _4744_ (.CLK(clk),
    .D(_0117_),
    .RESET_B(_0643_),
    .Q(out_data_flat[157]));
 sky130_fd_sc_hd__dfrtp_2 _4745_ (.CLK(clk),
    .D(_0119_),
    .RESET_B(_0644_),
    .Q(out_data_flat[158]));
 sky130_fd_sc_hd__dfrtp_2 _4746_ (.CLK(clk),
    .D(_0120_),
    .RESET_B(_0645_),
    .Q(out_data_flat[159]));
 sky130_fd_sc_hd__dfrtp_2 _4747_ (.CLK(clk),
    .D(_0064_),
    .RESET_B(_0646_),
    .Q(out_data_flat[96]));
 sky130_fd_sc_hd__dfrtp_2 _4748_ (.CLK(clk),
    .D(_0075_),
    .RESET_B(_0647_),
    .Q(out_data_flat[97]));
 sky130_fd_sc_hd__dfrtp_2 _4749_ (.CLK(clk),
    .D(_0086_),
    .RESET_B(_0648_),
    .Q(out_data_flat[98]));
 sky130_fd_sc_hd__dfrtp_2 _4750_ (.CLK(clk),
    .D(_0089_),
    .RESET_B(_0649_),
    .Q(out_data_flat[99]));
 sky130_fd_sc_hd__dfrtp_2 _4751_ (.CLK(clk),
    .D(_0090_),
    .RESET_B(_0650_),
    .Q(out_data_flat[100]));
 sky130_fd_sc_hd__dfrtp_2 _4752_ (.CLK(clk),
    .D(_0091_),
    .RESET_B(_0651_),
    .Q(out_data_flat[101]));
 sky130_fd_sc_hd__dfrtp_2 _4753_ (.CLK(clk),
    .D(_0092_),
    .RESET_B(_0652_),
    .Q(out_data_flat[102]));
 sky130_fd_sc_hd__dfrtp_2 _4754_ (.CLK(clk),
    .D(_0093_),
    .RESET_B(_0653_),
    .Q(out_data_flat[103]));
 sky130_fd_sc_hd__dfrtp_2 _4755_ (.CLK(clk),
    .D(_0094_),
    .RESET_B(_0654_),
    .Q(out_data_flat[104]));
 sky130_fd_sc_hd__dfrtp_2 _4756_ (.CLK(clk),
    .D(_0095_),
    .RESET_B(_0655_),
    .Q(out_data_flat[105]));
 sky130_fd_sc_hd__dfrtp_2 _4757_ (.CLK(clk),
    .D(_0065_),
    .RESET_B(_0656_),
    .Q(out_data_flat[106]));
 sky130_fd_sc_hd__dfrtp_2 _4758_ (.CLK(clk),
    .D(_0066_),
    .RESET_B(_0657_),
    .Q(out_data_flat[107]));
 sky130_fd_sc_hd__dfrtp_2 _4759_ (.CLK(clk),
    .D(_0067_),
    .RESET_B(_0658_),
    .Q(out_data_flat[108]));
 sky130_fd_sc_hd__dfrtp_2 _4760_ (.CLK(clk),
    .D(_0068_),
    .RESET_B(_0659_),
    .Q(out_data_flat[109]));
 sky130_fd_sc_hd__dfrtp_2 _4761_ (.CLK(clk),
    .D(_0069_),
    .RESET_B(_0660_),
    .Q(out_data_flat[110]));
 sky130_fd_sc_hd__dfrtp_2 _4762_ (.CLK(clk),
    .D(_0070_),
    .RESET_B(_0661_),
    .Q(out_data_flat[111]));
 sky130_fd_sc_hd__dfrtp_2 _4763_ (.CLK(clk),
    .D(_0071_),
    .RESET_B(_0662_),
    .Q(out_data_flat[112]));
 sky130_fd_sc_hd__dfrtp_2 _4764_ (.CLK(clk),
    .D(_0072_),
    .RESET_B(_0663_),
    .Q(out_data_flat[113]));
 sky130_fd_sc_hd__dfrtp_2 _4765_ (.CLK(clk),
    .D(_0073_),
    .RESET_B(_0664_),
    .Q(out_data_flat[114]));
 sky130_fd_sc_hd__dfrtp_2 _4766_ (.CLK(clk),
    .D(_0074_),
    .RESET_B(_0665_),
    .Q(out_data_flat[115]));
 sky130_fd_sc_hd__dfrtp_2 _4767_ (.CLK(clk),
    .D(_0076_),
    .RESET_B(_0666_),
    .Q(out_data_flat[116]));
 sky130_fd_sc_hd__dfrtp_2 _4768_ (.CLK(clk),
    .D(_0077_),
    .RESET_B(_0667_),
    .Q(out_data_flat[117]));
 sky130_fd_sc_hd__dfrtp_2 _4769_ (.CLK(clk),
    .D(_0078_),
    .RESET_B(_0668_),
    .Q(out_data_flat[118]));
 sky130_fd_sc_hd__dfrtp_2 _4770_ (.CLK(clk),
    .D(_0079_),
    .RESET_B(_0669_),
    .Q(out_data_flat[119]));
 sky130_fd_sc_hd__dfrtp_2 _4771_ (.CLK(clk),
    .D(_0080_),
    .RESET_B(_0670_),
    .Q(out_data_flat[120]));
 sky130_fd_sc_hd__dfrtp_2 _4772_ (.CLK(clk),
    .D(_0081_),
    .RESET_B(_0671_),
    .Q(out_data_flat[121]));
 sky130_fd_sc_hd__dfrtp_2 _4773_ (.CLK(clk),
    .D(_0082_),
    .RESET_B(_0672_),
    .Q(out_data_flat[122]));
 sky130_fd_sc_hd__dfrtp_2 _4774_ (.CLK(clk),
    .D(_0083_),
    .RESET_B(_0673_),
    .Q(out_data_flat[123]));
 sky130_fd_sc_hd__dfrtp_2 _4775_ (.CLK(clk),
    .D(_0084_),
    .RESET_B(_0674_),
    .Q(out_data_flat[124]));
 sky130_fd_sc_hd__dfrtp_2 _4776_ (.CLK(clk),
    .D(_0085_),
    .RESET_B(_0675_),
    .Q(out_data_flat[125]));
 sky130_fd_sc_hd__dfrtp_2 _4777_ (.CLK(clk),
    .D(_0087_),
    .RESET_B(_0676_),
    .Q(out_data_flat[126]));
 sky130_fd_sc_hd__dfrtp_2 _4778_ (.CLK(clk),
    .D(_0088_),
    .RESET_B(_0677_),
    .Q(out_data_flat[127]));
 sky130_fd_sc_hd__dfrtp_2 _4779_ (.CLK(clk),
    .D(_0032_),
    .RESET_B(_0678_),
    .Q(out_data_flat[64]));
 sky130_fd_sc_hd__dfrtp_2 _4780_ (.CLK(clk),
    .D(_0043_),
    .RESET_B(_0679_),
    .Q(out_data_flat[65]));
 sky130_fd_sc_hd__dfrtp_2 _4781_ (.CLK(clk),
    .D(_0054_),
    .RESET_B(_0680_),
    .Q(out_data_flat[66]));
 sky130_fd_sc_hd__dfrtp_2 _4782_ (.CLK(clk),
    .D(_0057_),
    .RESET_B(_0681_),
    .Q(out_data_flat[67]));
 sky130_fd_sc_hd__dfrtp_2 _4783_ (.CLK(clk),
    .D(_0058_),
    .RESET_B(_0682_),
    .Q(out_data_flat[68]));
 sky130_fd_sc_hd__dfrtp_2 _4784_ (.CLK(clk),
    .D(_0059_),
    .RESET_B(_0683_),
    .Q(out_data_flat[69]));
 sky130_fd_sc_hd__dfrtp_2 _4785_ (.CLK(clk),
    .D(_0060_),
    .RESET_B(_0684_),
    .Q(out_data_flat[70]));
 sky130_fd_sc_hd__dfrtp_2 _4786_ (.CLK(clk),
    .D(_0061_),
    .RESET_B(_0685_),
    .Q(out_data_flat[71]));
 sky130_fd_sc_hd__dfrtp_2 _4787_ (.CLK(clk),
    .D(_0062_),
    .RESET_B(_0686_),
    .Q(out_data_flat[72]));
 sky130_fd_sc_hd__dfrtp_2 _4788_ (.CLK(clk),
    .D(_0063_),
    .RESET_B(_0687_),
    .Q(out_data_flat[73]));
 sky130_fd_sc_hd__dfrtp_2 _4789_ (.CLK(clk),
    .D(_0033_),
    .RESET_B(_0688_),
    .Q(out_data_flat[74]));
 sky130_fd_sc_hd__dfrtp_2 _4790_ (.CLK(clk),
    .D(_0034_),
    .RESET_B(_0689_),
    .Q(out_data_flat[75]));
 sky130_fd_sc_hd__dfrtp_2 _4791_ (.CLK(clk),
    .D(_0035_),
    .RESET_B(_0690_),
    .Q(out_data_flat[76]));
 sky130_fd_sc_hd__dfrtp_2 _4792_ (.CLK(clk),
    .D(_0036_),
    .RESET_B(_0691_),
    .Q(out_data_flat[77]));
 sky130_fd_sc_hd__dfrtp_2 _4793_ (.CLK(clk),
    .D(_0037_),
    .RESET_B(_0692_),
    .Q(out_data_flat[78]));
 sky130_fd_sc_hd__dfrtp_2 _4794_ (.CLK(clk),
    .D(_0038_),
    .RESET_B(_0693_),
    .Q(out_data_flat[79]));
 sky130_fd_sc_hd__dfrtp_2 _4795_ (.CLK(clk),
    .D(_0039_),
    .RESET_B(_0694_),
    .Q(out_data_flat[80]));
 sky130_fd_sc_hd__dfrtp_2 _4796_ (.CLK(clk),
    .D(_0040_),
    .RESET_B(_0695_),
    .Q(out_data_flat[81]));
 sky130_fd_sc_hd__dfrtp_2 _4797_ (.CLK(clk),
    .D(_0041_),
    .RESET_B(_0696_),
    .Q(out_data_flat[82]));
 sky130_fd_sc_hd__dfrtp_2 _4798_ (.CLK(clk),
    .D(_0042_),
    .RESET_B(_0697_),
    .Q(out_data_flat[83]));
 sky130_fd_sc_hd__dfrtp_2 _4799_ (.CLK(clk),
    .D(_0044_),
    .RESET_B(_0698_),
    .Q(out_data_flat[84]));
 sky130_fd_sc_hd__dfrtp_2 _4800_ (.CLK(clk),
    .D(_0045_),
    .RESET_B(_0699_),
    .Q(out_data_flat[85]));
 sky130_fd_sc_hd__dfrtp_2 _4801_ (.CLK(clk),
    .D(_0046_),
    .RESET_B(_0700_),
    .Q(out_data_flat[86]));
 sky130_fd_sc_hd__dfrtp_2 _4802_ (.CLK(clk),
    .D(_0047_),
    .RESET_B(_0701_),
    .Q(out_data_flat[87]));
 sky130_fd_sc_hd__dfrtp_2 _4803_ (.CLK(clk),
    .D(_0048_),
    .RESET_B(_0702_),
    .Q(out_data_flat[88]));
 sky130_fd_sc_hd__dfrtp_2 _4804_ (.CLK(clk),
    .D(_0049_),
    .RESET_B(_0703_),
    .Q(out_data_flat[89]));
 sky130_fd_sc_hd__dfrtp_2 _4805_ (.CLK(clk),
    .D(_0050_),
    .RESET_B(_0704_),
    .Q(out_data_flat[90]));
 sky130_fd_sc_hd__dfrtp_2 _4806_ (.CLK(clk),
    .D(_0051_),
    .RESET_B(_0705_),
    .Q(out_data_flat[91]));
 sky130_fd_sc_hd__dfrtp_2 _4807_ (.CLK(clk),
    .D(_0052_),
    .RESET_B(_0706_),
    .Q(out_data_flat[92]));
 sky130_fd_sc_hd__dfrtp_2 _4808_ (.CLK(clk),
    .D(_0053_),
    .RESET_B(_0707_),
    .Q(out_data_flat[93]));
 sky130_fd_sc_hd__dfrtp_2 _4809_ (.CLK(clk),
    .D(_0055_),
    .RESET_B(_0708_),
    .Q(out_data_flat[94]));
 sky130_fd_sc_hd__dfrtp_2 _4810_ (.CLK(clk),
    .D(_0056_),
    .RESET_B(_0709_),
    .Q(out_data_flat[95]));
 sky130_fd_sc_hd__dfrtp_2 _4811_ (.CLK(clk),
    .D(_0000_),
    .RESET_B(_0710_),
    .Q(out_data_flat[32]));
 sky130_fd_sc_hd__dfrtp_2 _4812_ (.CLK(clk),
    .D(_0011_),
    .RESET_B(_0711_),
    .Q(out_data_flat[33]));
 sky130_fd_sc_hd__dfrtp_2 _4813_ (.CLK(clk),
    .D(_0022_),
    .RESET_B(_0712_),
    .Q(out_data_flat[34]));
 sky130_fd_sc_hd__dfrtp_2 _4814_ (.CLK(clk),
    .D(_0025_),
    .RESET_B(_0713_),
    .Q(out_data_flat[35]));
 sky130_fd_sc_hd__dfrtp_2 _4815_ (.CLK(clk),
    .D(_0026_),
    .RESET_B(_0714_),
    .Q(out_data_flat[36]));
 sky130_fd_sc_hd__dfrtp_2 _4816_ (.CLK(clk),
    .D(_0027_),
    .RESET_B(_0715_),
    .Q(out_data_flat[37]));
 sky130_fd_sc_hd__dfrtp_2 _4817_ (.CLK(clk),
    .D(_0028_),
    .RESET_B(_0716_),
    .Q(out_data_flat[38]));
 sky130_fd_sc_hd__dfrtp_2 _4818_ (.CLK(clk),
    .D(_0029_),
    .RESET_B(_0717_),
    .Q(out_data_flat[39]));
 sky130_fd_sc_hd__dfrtp_2 _4819_ (.CLK(clk),
    .D(_0030_),
    .RESET_B(_0718_),
    .Q(out_data_flat[40]));
 sky130_fd_sc_hd__dfrtp_2 _4820_ (.CLK(clk),
    .D(_0031_),
    .RESET_B(_0719_),
    .Q(out_data_flat[41]));
 sky130_fd_sc_hd__dfrtp_2 _4821_ (.CLK(clk),
    .D(_0001_),
    .RESET_B(_0720_),
    .Q(out_data_flat[42]));
 sky130_fd_sc_hd__dfrtp_2 _4822_ (.CLK(clk),
    .D(_0002_),
    .RESET_B(_0721_),
    .Q(out_data_flat[43]));
 sky130_fd_sc_hd__dfrtp_2 _4823_ (.CLK(clk),
    .D(_0003_),
    .RESET_B(_0722_),
    .Q(out_data_flat[44]));
 sky130_fd_sc_hd__dfrtp_2 _4824_ (.CLK(clk),
    .D(_0004_),
    .RESET_B(_0723_),
    .Q(out_data_flat[45]));
 sky130_fd_sc_hd__dfrtp_2 _4825_ (.CLK(clk),
    .D(_0005_),
    .RESET_B(_0724_),
    .Q(out_data_flat[46]));
 sky130_fd_sc_hd__dfrtp_2 _4826_ (.CLK(clk),
    .D(_0006_),
    .RESET_B(_0725_),
    .Q(out_data_flat[47]));
 sky130_fd_sc_hd__dfrtp_2 _4827_ (.CLK(clk),
    .D(_0007_),
    .RESET_B(_0726_),
    .Q(out_data_flat[48]));
 sky130_fd_sc_hd__dfrtp_2 _4828_ (.CLK(clk),
    .D(_0008_),
    .RESET_B(_0727_),
    .Q(out_data_flat[49]));
 sky130_fd_sc_hd__dfrtp_2 _4829_ (.CLK(clk),
    .D(_0009_),
    .RESET_B(_0728_),
    .Q(out_data_flat[50]));
 sky130_fd_sc_hd__dfrtp_2 _4830_ (.CLK(clk),
    .D(_0010_),
    .RESET_B(_0729_),
    .Q(out_data_flat[51]));
 sky130_fd_sc_hd__dfrtp_2 _4831_ (.CLK(clk),
    .D(_0012_),
    .RESET_B(_0730_),
    .Q(out_data_flat[52]));
 sky130_fd_sc_hd__dfrtp_2 _4832_ (.CLK(clk),
    .D(_0013_),
    .RESET_B(_0731_),
    .Q(out_data_flat[53]));
 sky130_fd_sc_hd__dfrtp_2 _4833_ (.CLK(clk),
    .D(_0014_),
    .RESET_B(_0732_),
    .Q(out_data_flat[54]));
 sky130_fd_sc_hd__dfrtp_2 _4834_ (.CLK(clk),
    .D(_0015_),
    .RESET_B(_0733_),
    .Q(out_data_flat[55]));
 sky130_fd_sc_hd__dfrtp_2 _4835_ (.CLK(clk),
    .D(_0016_),
    .RESET_B(_0734_),
    .Q(out_data_flat[56]));
 sky130_fd_sc_hd__dfrtp_2 _4836_ (.CLK(clk),
    .D(_0017_),
    .RESET_B(_0735_),
    .Q(out_data_flat[57]));
 sky130_fd_sc_hd__dfrtp_2 _4837_ (.CLK(clk),
    .D(_0018_),
    .RESET_B(_0736_),
    .Q(out_data_flat[58]));
 sky130_fd_sc_hd__dfrtp_2 _4838_ (.CLK(clk),
    .D(_0019_),
    .RESET_B(_0737_),
    .Q(out_data_flat[59]));
 sky130_fd_sc_hd__dfrtp_2 _4839_ (.CLK(clk),
    .D(_0020_),
    .RESET_B(_0738_),
    .Q(out_data_flat[60]));
 sky130_fd_sc_hd__dfrtp_2 _4840_ (.CLK(clk),
    .D(_0021_),
    .RESET_B(_0739_),
    .Q(out_data_flat[61]));
 sky130_fd_sc_hd__dfrtp_2 _4841_ (.CLK(clk),
    .D(_0023_),
    .RESET_B(_0740_),
    .Q(out_data_flat[62]));
 sky130_fd_sc_hd__dfrtp_2 _4842_ (.CLK(clk),
    .D(_0024_),
    .RESET_B(_0741_),
    .Q(out_data_flat[63]));
 sky130_fd_sc_hd__dfrtp_2 _4843_ (.CLK(clk),
    .D(_0192_),
    .RESET_B(_0742_),
    .Q(\gen_pe[1].pe_inst.sel ));
 sky130_fd_sc_hd__dfrtp_2 _4844_ (.CLK(clk),
    .D(_0609_),
    .RESET_B(_0743_),
    .Q(\gen_pe[6].pe_inst.out_right[0] ));
 sky130_fd_sc_hd__dfrtp_2 _4845_ (.CLK(clk),
    .D(_0620_),
    .RESET_B(_0744_),
    .Q(\gen_pe[6].pe_inst.out_right[1] ));
 sky130_fd_sc_hd__dfrtp_2 _4846_ (.CLK(clk),
    .D(_0631_),
    .RESET_B(_0745_),
    .Q(\gen_pe[6].pe_inst.out_right[2] ));
 sky130_fd_sc_hd__dfrtp_2 _4847_ (.CLK(clk),
    .D(_0634_),
    .RESET_B(_0746_),
    .Q(\gen_pe[6].pe_inst.out_right[3] ));
 sky130_fd_sc_hd__dfrtp_2 _4848_ (.CLK(clk),
    .D(_0635_),
    .RESET_B(_0747_),
    .Q(\gen_pe[6].pe_inst.out_right[4] ));
 sky130_fd_sc_hd__dfrtp_2 _4849_ (.CLK(clk),
    .D(_0636_),
    .RESET_B(_0748_),
    .Q(\gen_pe[6].pe_inst.out_right[5] ));
 sky130_fd_sc_hd__dfrtp_2 _4850_ (.CLK(clk),
    .D(_0637_),
    .RESET_B(_0749_),
    .Q(\gen_pe[6].pe_inst.out_right[6] ));
 sky130_fd_sc_hd__dfrtp_2 _4851_ (.CLK(clk),
    .D(_0638_),
    .RESET_B(_0750_),
    .Q(\gen_pe[6].pe_inst.out_right[7] ));
 sky130_fd_sc_hd__dfrtp_2 _4852_ (.CLK(clk),
    .D(_0639_),
    .RESET_B(_0751_),
    .Q(\gen_pe[6].pe_inst.out_right[8] ));
 sky130_fd_sc_hd__dfrtp_2 _4853_ (.CLK(clk),
    .D(_0640_),
    .RESET_B(_0752_),
    .Q(\gen_pe[6].pe_inst.out_right[9] ));
 sky130_fd_sc_hd__dfrtp_2 _4854_ (.CLK(clk),
    .D(_0610_),
    .RESET_B(_0753_),
    .Q(\gen_pe[6].pe_inst.out_right[10] ));
 sky130_fd_sc_hd__dfrtp_2 _4855_ (.CLK(clk),
    .D(_0611_),
    .RESET_B(_0754_),
    .Q(\gen_pe[6].pe_inst.out_right[11] ));
 sky130_fd_sc_hd__dfrtp_2 _4856_ (.CLK(clk),
    .D(_0612_),
    .RESET_B(_0755_),
    .Q(\gen_pe[6].pe_inst.out_right[12] ));
 sky130_fd_sc_hd__dfrtp_2 _4857_ (.CLK(clk),
    .D(_0613_),
    .RESET_B(_0756_),
    .Q(\gen_pe[6].pe_inst.out_right[13] ));
 sky130_fd_sc_hd__dfrtp_2 _4858_ (.CLK(clk),
    .D(_0614_),
    .RESET_B(_0757_),
    .Q(\gen_pe[6].pe_inst.out_right[14] ));
 sky130_fd_sc_hd__dfrtp_2 _4859_ (.CLK(clk),
    .D(_0615_),
    .RESET_B(_0758_),
    .Q(\gen_pe[6].pe_inst.out_right[15] ));
 sky130_fd_sc_hd__dfrtp_2 _4860_ (.CLK(clk),
    .D(_0616_),
    .RESET_B(_0759_),
    .Q(\gen_pe[6].pe_inst.out_right[16] ));
 sky130_fd_sc_hd__dfrtp_2 _4861_ (.CLK(clk),
    .D(_0617_),
    .RESET_B(_0760_),
    .Q(\gen_pe[6].pe_inst.out_right[17] ));
 sky130_fd_sc_hd__dfrtp_2 _4862_ (.CLK(clk),
    .D(_0618_),
    .RESET_B(_0761_),
    .Q(\gen_pe[6].pe_inst.out_right[18] ));
 sky130_fd_sc_hd__dfrtp_2 _4863_ (.CLK(clk),
    .D(_0619_),
    .RESET_B(_0762_),
    .Q(\gen_pe[6].pe_inst.out_right[19] ));
 sky130_fd_sc_hd__dfrtp_2 _4864_ (.CLK(clk),
    .D(_0621_),
    .RESET_B(_0763_),
    .Q(\gen_pe[6].pe_inst.out_right[20] ));
 sky130_fd_sc_hd__dfrtp_2 _4865_ (.CLK(clk),
    .D(_0622_),
    .RESET_B(_0764_),
    .Q(\gen_pe[6].pe_inst.out_right[21] ));
 sky130_fd_sc_hd__dfrtp_2 _4866_ (.CLK(clk),
    .D(_0623_),
    .RESET_B(_0765_),
    .Q(\gen_pe[6].pe_inst.out_right[22] ));
 sky130_fd_sc_hd__dfrtp_2 _4867_ (.CLK(clk),
    .D(_0624_),
    .RESET_B(_0766_),
    .Q(\gen_pe[6].pe_inst.out_right[23] ));
 sky130_fd_sc_hd__dfrtp_2 _4868_ (.CLK(clk),
    .D(_0625_),
    .RESET_B(_0767_),
    .Q(\gen_pe[6].pe_inst.out_right[24] ));
 sky130_fd_sc_hd__dfrtp_2 _4869_ (.CLK(clk),
    .D(_0626_),
    .RESET_B(_0768_),
    .Q(\gen_pe[6].pe_inst.out_right[25] ));
 sky130_fd_sc_hd__dfrtp_2 _4870_ (.CLK(clk),
    .D(_0627_),
    .RESET_B(_0769_),
    .Q(\gen_pe[6].pe_inst.out_right[26] ));
 sky130_fd_sc_hd__dfrtp_2 _4871_ (.CLK(clk),
    .D(_0628_),
    .RESET_B(_0770_),
    .Q(\gen_pe[6].pe_inst.out_right[27] ));
 sky130_fd_sc_hd__dfrtp_2 _4872_ (.CLK(clk),
    .D(_0629_),
    .RESET_B(_0771_),
    .Q(\gen_pe[6].pe_inst.out_right[28] ));
 sky130_fd_sc_hd__dfrtp_2 _4873_ (.CLK(clk),
    .D(_0630_),
    .RESET_B(_0772_),
    .Q(\gen_pe[6].pe_inst.out_right[29] ));
 sky130_fd_sc_hd__dfrtp_2 _4874_ (.CLK(clk),
    .D(_0632_),
    .RESET_B(_0773_),
    .Q(\gen_pe[6].pe_inst.out_right[30] ));
 sky130_fd_sc_hd__dfrtp_2 _4875_ (.CLK(clk),
    .D(_0633_),
    .RESET_B(_0774_),
    .Q(\gen_pe[6].pe_inst.out_right[31] ));
 sky130_fd_sc_hd__dfrtp_2 _4876_ (.CLK(clk),
    .D(_0289_),
    .RESET_B(_0775_),
    .Q(\gen_pe[1].pe_inst.out_right[0] ));
 sky130_fd_sc_hd__dfrtp_2 _4877_ (.CLK(clk),
    .D(_0300_),
    .RESET_B(_0776_),
    .Q(\gen_pe[1].pe_inst.out_right[1] ));
 sky130_fd_sc_hd__dfrtp_2 _4878_ (.CLK(clk),
    .D(_0311_),
    .RESET_B(_0777_),
    .Q(\gen_pe[1].pe_inst.out_right[2] ));
 sky130_fd_sc_hd__dfrtp_2 _4879_ (.CLK(clk),
    .D(_0314_),
    .RESET_B(_0778_),
    .Q(\gen_pe[1].pe_inst.out_right[3] ));
 sky130_fd_sc_hd__dfrtp_2 _4880_ (.CLK(clk),
    .D(_0315_),
    .RESET_B(_0779_),
    .Q(\gen_pe[1].pe_inst.out_right[4] ));
 sky130_fd_sc_hd__dfrtp_2 _4881_ (.CLK(clk),
    .D(_0316_),
    .RESET_B(_0780_),
    .Q(\gen_pe[1].pe_inst.out_right[5] ));
 sky130_fd_sc_hd__dfrtp_2 _4882_ (.CLK(clk),
    .D(_0317_),
    .RESET_B(_0781_),
    .Q(\gen_pe[1].pe_inst.out_right[6] ));
 sky130_fd_sc_hd__dfrtp_2 _4883_ (.CLK(clk),
    .D(_0318_),
    .RESET_B(_0782_),
    .Q(\gen_pe[1].pe_inst.out_right[7] ));
 sky130_fd_sc_hd__dfrtp_2 _4884_ (.CLK(clk),
    .D(_0319_),
    .RESET_B(_0783_),
    .Q(\gen_pe[1].pe_inst.out_right[8] ));
 sky130_fd_sc_hd__dfrtp_2 _4885_ (.CLK(clk),
    .D(_0320_),
    .RESET_B(_0784_),
    .Q(\gen_pe[1].pe_inst.out_right[9] ));
 sky130_fd_sc_hd__dfrtp_2 _4886_ (.CLK(clk),
    .D(_0290_),
    .RESET_B(_0785_),
    .Q(\gen_pe[1].pe_inst.out_right[10] ));
 sky130_fd_sc_hd__dfrtp_2 _4887_ (.CLK(clk),
    .D(_0291_),
    .RESET_B(_0786_),
    .Q(\gen_pe[1].pe_inst.out_right[11] ));
 sky130_fd_sc_hd__dfrtp_2 _4888_ (.CLK(clk),
    .D(_0292_),
    .RESET_B(_0787_),
    .Q(\gen_pe[1].pe_inst.out_right[12] ));
 sky130_fd_sc_hd__dfrtp_2 _4889_ (.CLK(clk),
    .D(_0293_),
    .RESET_B(_0788_),
    .Q(\gen_pe[1].pe_inst.out_right[13] ));
 sky130_fd_sc_hd__dfrtp_2 _4890_ (.CLK(clk),
    .D(_0294_),
    .RESET_B(_0789_),
    .Q(\gen_pe[1].pe_inst.out_right[14] ));
 sky130_fd_sc_hd__dfrtp_2 _4891_ (.CLK(clk),
    .D(_0295_),
    .RESET_B(_0790_),
    .Q(\gen_pe[1].pe_inst.out_right[15] ));
 sky130_fd_sc_hd__dfrtp_2 _4892_ (.CLK(clk),
    .D(_0296_),
    .RESET_B(_0791_),
    .Q(\gen_pe[1].pe_inst.out_right[16] ));
 sky130_fd_sc_hd__dfrtp_2 _4893_ (.CLK(clk),
    .D(_0297_),
    .RESET_B(_0792_),
    .Q(\gen_pe[1].pe_inst.out_right[17] ));
 sky130_fd_sc_hd__dfrtp_2 _4894_ (.CLK(clk),
    .D(_0298_),
    .RESET_B(_0793_),
    .Q(\gen_pe[1].pe_inst.out_right[18] ));
 sky130_fd_sc_hd__dfrtp_2 _4895_ (.CLK(clk),
    .D(_0299_),
    .RESET_B(_0794_),
    .Q(\gen_pe[1].pe_inst.out_right[19] ));
 sky130_fd_sc_hd__dfrtp_2 _4896_ (.CLK(clk),
    .D(_0301_),
    .RESET_B(_0795_),
    .Q(\gen_pe[1].pe_inst.out_right[20] ));
 sky130_fd_sc_hd__dfrtp_2 _4897_ (.CLK(clk),
    .D(_0302_),
    .RESET_B(_0796_),
    .Q(\gen_pe[1].pe_inst.out_right[21] ));
 sky130_fd_sc_hd__dfrtp_2 _4898_ (.CLK(clk),
    .D(_0303_),
    .RESET_B(_0797_),
    .Q(\gen_pe[1].pe_inst.out_right[22] ));
 sky130_fd_sc_hd__dfrtp_2 _4899_ (.CLK(clk),
    .D(_0304_),
    .RESET_B(_0798_),
    .Q(\gen_pe[1].pe_inst.out_right[23] ));
 sky130_fd_sc_hd__dfrtp_2 _4900_ (.CLK(clk),
    .D(_0305_),
    .RESET_B(_0799_),
    .Q(\gen_pe[1].pe_inst.out_right[24] ));
 sky130_fd_sc_hd__dfrtp_2 _4901_ (.CLK(clk),
    .D(_0306_),
    .RESET_B(_0800_),
    .Q(\gen_pe[1].pe_inst.out_right[25] ));
 sky130_fd_sc_hd__dfrtp_2 _4902_ (.CLK(clk),
    .D(_0307_),
    .RESET_B(_0801_),
    .Q(\gen_pe[1].pe_inst.out_right[26] ));
 sky130_fd_sc_hd__dfrtp_2 _4903_ (.CLK(clk),
    .D(_0308_),
    .RESET_B(_0802_),
    .Q(\gen_pe[1].pe_inst.out_right[27] ));
 sky130_fd_sc_hd__dfrtp_2 _4904_ (.CLK(clk),
    .D(_0309_),
    .RESET_B(_0803_),
    .Q(\gen_pe[1].pe_inst.out_right[28] ));
 sky130_fd_sc_hd__dfrtp_2 _4905_ (.CLK(clk),
    .D(_0310_),
    .RESET_B(_0804_),
    .Q(\gen_pe[1].pe_inst.out_right[29] ));
 sky130_fd_sc_hd__dfrtp_2 _4906_ (.CLK(clk),
    .D(_0312_),
    .RESET_B(_0805_),
    .Q(\gen_pe[1].pe_inst.out_right[30] ));
 sky130_fd_sc_hd__dfrtp_2 _4907_ (.CLK(clk),
    .D(_0313_),
    .RESET_B(_0806_),
    .Q(\gen_pe[1].pe_inst.out_right[31] ));
 sky130_fd_sc_hd__dfrtp_2 _4908_ (.CLK(clk),
    .D(_0257_),
    .RESET_B(_0807_),
    .Q(\gen_left[1][0] ));
 sky130_fd_sc_hd__dfrtp_2 _4909_ (.CLK(clk),
    .D(_0268_),
    .RESET_B(_0808_),
    .Q(\gen_left[1][1] ));
 sky130_fd_sc_hd__dfrtp_2 _4910_ (.CLK(clk),
    .D(_0279_),
    .RESET_B(_0809_),
    .Q(\gen_left[1][2] ));
 sky130_fd_sc_hd__dfrtp_2 _4911_ (.CLK(clk),
    .D(_0282_),
    .RESET_B(_0810_),
    .Q(\gen_left[1][3] ));
 sky130_fd_sc_hd__dfrtp_2 _4912_ (.CLK(clk),
    .D(_0283_),
    .RESET_B(_0811_),
    .Q(\gen_left[1][4] ));
 sky130_fd_sc_hd__dfrtp_2 _4913_ (.CLK(clk),
    .D(_0284_),
    .RESET_B(_0812_),
    .Q(\gen_left[1][5] ));
 sky130_fd_sc_hd__dfrtp_2 _4914_ (.CLK(clk),
    .D(_0285_),
    .RESET_B(_0813_),
    .Q(\gen_left[1][6] ));
 sky130_fd_sc_hd__dfrtp_2 _4915_ (.CLK(clk),
    .D(_0286_),
    .RESET_B(_0814_),
    .Q(\gen_left[1][7] ));
 sky130_fd_sc_hd__dfrtp_2 _4916_ (.CLK(clk),
    .D(_0287_),
    .RESET_B(_0815_),
    .Q(\gen_left[1][8] ));
 sky130_fd_sc_hd__dfrtp_2 _4917_ (.CLK(clk),
    .D(_0288_),
    .RESET_B(_0816_),
    .Q(\gen_left[1][9] ));
 sky130_fd_sc_hd__dfrtp_2 _4918_ (.CLK(clk),
    .D(_0258_),
    .RESET_B(_0817_),
    .Q(\gen_left[1][10] ));
 sky130_fd_sc_hd__dfrtp_2 _4919_ (.CLK(clk),
    .D(_0259_),
    .RESET_B(_0818_),
    .Q(\gen_left[1][11] ));
 sky130_fd_sc_hd__dfrtp_2 _4920_ (.CLK(clk),
    .D(_0260_),
    .RESET_B(_0819_),
    .Q(\gen_left[1][12] ));
 sky130_fd_sc_hd__dfrtp_2 _4921_ (.CLK(clk),
    .D(_0261_),
    .RESET_B(_0820_),
    .Q(\gen_left[1][13] ));
 sky130_fd_sc_hd__dfrtp_2 _4922_ (.CLK(clk),
    .D(_0262_),
    .RESET_B(_0821_),
    .Q(\gen_left[1][14] ));
 sky130_fd_sc_hd__dfrtp_2 _4923_ (.CLK(clk),
    .D(_0263_),
    .RESET_B(_0822_),
    .Q(\gen_left[1][15] ));
 sky130_fd_sc_hd__dfrtp_2 _4924_ (.CLK(clk),
    .D(_0264_),
    .RESET_B(_0823_),
    .Q(\gen_left[1][16] ));
 sky130_fd_sc_hd__dfrtp_2 _4925_ (.CLK(clk),
    .D(_0265_),
    .RESET_B(_0824_),
    .Q(\gen_left[1][17] ));
 sky130_fd_sc_hd__dfrtp_2 _4926_ (.CLK(clk),
    .D(_0266_),
    .RESET_B(_0825_),
    .Q(\gen_left[1][18] ));
 sky130_fd_sc_hd__dfrtp_2 _4927_ (.CLK(clk),
    .D(_0267_),
    .RESET_B(_0826_),
    .Q(\gen_left[1][19] ));
 sky130_fd_sc_hd__dfrtp_2 _4928_ (.CLK(clk),
    .D(_0269_),
    .RESET_B(_0827_),
    .Q(\gen_left[1][20] ));
 sky130_fd_sc_hd__dfrtp_2 _4929_ (.CLK(clk),
    .D(_0270_),
    .RESET_B(_0828_),
    .Q(\gen_left[1][21] ));
 sky130_fd_sc_hd__dfrtp_2 _4930_ (.CLK(clk),
    .D(_0271_),
    .RESET_B(_0829_),
    .Q(\gen_left[1][22] ));
 sky130_fd_sc_hd__dfrtp_2 _4931_ (.CLK(clk),
    .D(_0272_),
    .RESET_B(_0830_),
    .Q(\gen_left[1][23] ));
 sky130_fd_sc_hd__dfrtp_2 _4932_ (.CLK(clk),
    .D(_0273_),
    .RESET_B(_0831_),
    .Q(\gen_left[1][24] ));
 sky130_fd_sc_hd__dfrtp_2 _4933_ (.CLK(clk),
    .D(_0274_),
    .RESET_B(_0832_),
    .Q(\gen_left[1][25] ));
 sky130_fd_sc_hd__dfrtp_2 _4934_ (.CLK(clk),
    .D(_0275_),
    .RESET_B(_0833_),
    .Q(\gen_left[1][26] ));
 sky130_fd_sc_hd__dfrtp_2 _4935_ (.CLK(clk),
    .D(_0276_),
    .RESET_B(_0834_),
    .Q(\gen_left[1][27] ));
 sky130_fd_sc_hd__dfrtp_2 _4936_ (.CLK(clk),
    .D(_0277_),
    .RESET_B(_0835_),
    .Q(\gen_left[1][28] ));
 sky130_fd_sc_hd__dfrtp_2 _4937_ (.CLK(clk),
    .D(_0278_),
    .RESET_B(_0836_),
    .Q(\gen_left[1][29] ));
 sky130_fd_sc_hd__dfrtp_2 _4938_ (.CLK(clk),
    .D(_0280_),
    .RESET_B(_0837_),
    .Q(\gen_left[1][30] ));
 sky130_fd_sc_hd__dfrtp_2 _4939_ (.CLK(clk),
    .D(_0281_),
    .RESET_B(_0838_),
    .Q(\gen_left[1][31] ));
 sky130_fd_sc_hd__dfrtp_2 _4940_ (.CLK(clk),
    .D(_0225_),
    .RESET_B(_0839_),
    .Q(\gen_pe[0].pe_inst.out_right[0] ));
 sky130_fd_sc_hd__dfrtp_2 _4941_ (.CLK(clk),
    .D(_0236_),
    .RESET_B(_0840_),
    .Q(\gen_pe[0].pe_inst.out_right[1] ));
 sky130_fd_sc_hd__dfrtp_2 _4942_ (.CLK(clk),
    .D(_0247_),
    .RESET_B(_0841_),
    .Q(\gen_pe[0].pe_inst.out_right[2] ));
 sky130_fd_sc_hd__dfrtp_2 _4943_ (.CLK(clk),
    .D(_0250_),
    .RESET_B(_0842_),
    .Q(\gen_pe[0].pe_inst.out_right[3] ));
 sky130_fd_sc_hd__dfrtp_2 _4944_ (.CLK(clk),
    .D(_0251_),
    .RESET_B(_0843_),
    .Q(\gen_pe[0].pe_inst.out_right[4] ));
 sky130_fd_sc_hd__dfrtp_2 _4945_ (.CLK(clk),
    .D(_0252_),
    .RESET_B(_0844_),
    .Q(\gen_pe[0].pe_inst.out_right[5] ));
 sky130_fd_sc_hd__dfrtp_2 _4946_ (.CLK(clk),
    .D(_0253_),
    .RESET_B(_0845_),
    .Q(\gen_pe[0].pe_inst.out_right[6] ));
 sky130_fd_sc_hd__dfrtp_2 _4947_ (.CLK(clk),
    .D(_0254_),
    .RESET_B(_0846_),
    .Q(\gen_pe[0].pe_inst.out_right[7] ));
 sky130_fd_sc_hd__dfrtp_2 _4948_ (.CLK(clk),
    .D(_0255_),
    .RESET_B(_0847_),
    .Q(\gen_pe[0].pe_inst.out_right[8] ));
 sky130_fd_sc_hd__dfrtp_2 _4949_ (.CLK(clk),
    .D(_0256_),
    .RESET_B(_0848_),
    .Q(\gen_pe[0].pe_inst.out_right[9] ));
 sky130_fd_sc_hd__dfrtp_2 _4950_ (.CLK(clk),
    .D(_0226_),
    .RESET_B(_0849_),
    .Q(\gen_pe[0].pe_inst.out_right[10] ));
 sky130_fd_sc_hd__dfrtp_2 _4951_ (.CLK(clk),
    .D(_0227_),
    .RESET_B(_0850_),
    .Q(\gen_pe[0].pe_inst.out_right[11] ));
 sky130_fd_sc_hd__dfrtp_2 _4952_ (.CLK(clk),
    .D(_0228_),
    .RESET_B(_0851_),
    .Q(\gen_pe[0].pe_inst.out_right[12] ));
 sky130_fd_sc_hd__dfrtp_2 _4953_ (.CLK(clk),
    .D(_0229_),
    .RESET_B(_0852_),
    .Q(\gen_pe[0].pe_inst.out_right[13] ));
 sky130_fd_sc_hd__dfrtp_2 _4954_ (.CLK(clk),
    .D(_0230_),
    .RESET_B(_0853_),
    .Q(\gen_pe[0].pe_inst.out_right[14] ));
 sky130_fd_sc_hd__dfrtp_2 _4955_ (.CLK(clk),
    .D(_0231_),
    .RESET_B(_0854_),
    .Q(\gen_pe[0].pe_inst.out_right[15] ));
 sky130_fd_sc_hd__dfrtp_2 _4956_ (.CLK(clk),
    .D(_0232_),
    .RESET_B(_0855_),
    .Q(\gen_pe[0].pe_inst.out_right[16] ));
 sky130_fd_sc_hd__dfrtp_2 _4957_ (.CLK(clk),
    .D(_0233_),
    .RESET_B(_0856_),
    .Q(\gen_pe[0].pe_inst.out_right[17] ));
 sky130_fd_sc_hd__dfrtp_2 _4958_ (.CLK(clk),
    .D(_0234_),
    .RESET_B(_0857_),
    .Q(\gen_pe[0].pe_inst.out_right[18] ));
 sky130_fd_sc_hd__dfrtp_2 _4959_ (.CLK(clk),
    .D(_0235_),
    .RESET_B(_0858_),
    .Q(\gen_pe[0].pe_inst.out_right[19] ));
 sky130_fd_sc_hd__dfrtp_2 _4960_ (.CLK(clk),
    .D(_0237_),
    .RESET_B(_0859_),
    .Q(\gen_pe[0].pe_inst.out_right[20] ));
 sky130_fd_sc_hd__dfrtp_2 _4961_ (.CLK(clk),
    .D(_0238_),
    .RESET_B(_0860_),
    .Q(\gen_pe[0].pe_inst.out_right[21] ));
 sky130_fd_sc_hd__dfrtp_2 _4962_ (.CLK(clk),
    .D(_0239_),
    .RESET_B(_0861_),
    .Q(\gen_pe[0].pe_inst.out_right[22] ));
 sky130_fd_sc_hd__dfrtp_2 _4963_ (.CLK(clk),
    .D(_0240_),
    .RESET_B(_0862_),
    .Q(\gen_pe[0].pe_inst.out_right[23] ));
 sky130_fd_sc_hd__dfrtp_2 _4964_ (.CLK(clk),
    .D(_0241_),
    .RESET_B(_0863_),
    .Q(\gen_pe[0].pe_inst.out_right[24] ));
 sky130_fd_sc_hd__dfrtp_2 _4965_ (.CLK(clk),
    .D(_0242_),
    .RESET_B(_0864_),
    .Q(\gen_pe[0].pe_inst.out_right[25] ));
 sky130_fd_sc_hd__dfrtp_2 _4966_ (.CLK(clk),
    .D(_0243_),
    .RESET_B(_0865_),
    .Q(\gen_pe[0].pe_inst.out_right[26] ));
 sky130_fd_sc_hd__dfrtp_2 _4967_ (.CLK(clk),
    .D(_0244_),
    .RESET_B(_0866_),
    .Q(\gen_pe[0].pe_inst.out_right[27] ));
 sky130_fd_sc_hd__dfrtp_2 _4968_ (.CLK(clk),
    .D(_0245_),
    .RESET_B(_0867_),
    .Q(\gen_pe[0].pe_inst.out_right[28] ));
 sky130_fd_sc_hd__dfrtp_2 _4969_ (.CLK(clk),
    .D(_0246_),
    .RESET_B(_0868_),
    .Q(\gen_pe[0].pe_inst.out_right[29] ));
 sky130_fd_sc_hd__dfrtp_2 _4970_ (.CLK(clk),
    .D(_0248_),
    .RESET_B(_0869_),
    .Q(\gen_pe[0].pe_inst.out_right[30] ));
 sky130_fd_sc_hd__dfrtp_2 _4971_ (.CLK(clk),
    .D(_0249_),
    .RESET_B(_0870_),
    .Q(\gen_pe[0].pe_inst.out_right[31] ));
 sky130_fd_sc_hd__dfrtp_2 _4972_ (.CLK(clk),
    .D(_0193_),
    .RESET_B(_0871_),
    .Q(\gen_left[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _4973_ (.CLK(clk),
    .D(_0204_),
    .RESET_B(_0872_),
    .Q(\gen_left[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _4974_ (.CLK(clk),
    .D(_0215_),
    .RESET_B(_0873_),
    .Q(\gen_left[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _4975_ (.CLK(clk),
    .D(_0218_),
    .RESET_B(_0874_),
    .Q(\gen_left[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _4976_ (.CLK(clk),
    .D(_0219_),
    .RESET_B(_0875_),
    .Q(\gen_left[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _4977_ (.CLK(clk),
    .D(_0220_),
    .RESET_B(_0876_),
    .Q(\gen_left[0][5] ));
 sky130_fd_sc_hd__dfrtp_2 _4978_ (.CLK(clk),
    .D(_0221_),
    .RESET_B(_0877_),
    .Q(\gen_left[0][6] ));
 sky130_fd_sc_hd__dfrtp_2 _4979_ (.CLK(clk),
    .D(_0222_),
    .RESET_B(_0878_),
    .Q(\gen_left[0][7] ));
 sky130_fd_sc_hd__dfrtp_2 _4980_ (.CLK(clk),
    .D(_0223_),
    .RESET_B(_0879_),
    .Q(\gen_left[0][8] ));
 sky130_fd_sc_hd__dfrtp_2 _4981_ (.CLK(clk),
    .D(_0224_),
    .RESET_B(_0880_),
    .Q(\gen_left[0][9] ));
 sky130_fd_sc_hd__dfrtp_2 _4982_ (.CLK(clk),
    .D(_0194_),
    .RESET_B(_0881_),
    .Q(\gen_left[0][10] ));
 sky130_fd_sc_hd__dfrtp_2 _4983_ (.CLK(clk),
    .D(_0195_),
    .RESET_B(_0882_),
    .Q(\gen_left[0][11] ));
 sky130_fd_sc_hd__dfrtp_2 _4984_ (.CLK(clk),
    .D(_0196_),
    .RESET_B(_0883_),
    .Q(\gen_left[0][12] ));
 sky130_fd_sc_hd__dfrtp_2 _4985_ (.CLK(clk),
    .D(_0197_),
    .RESET_B(_0884_),
    .Q(\gen_left[0][13] ));
 sky130_fd_sc_hd__dfrtp_2 _4986_ (.CLK(clk),
    .D(_0198_),
    .RESET_B(_0885_),
    .Q(\gen_left[0][14] ));
 sky130_fd_sc_hd__dfrtp_2 _4987_ (.CLK(clk),
    .D(_0199_),
    .RESET_B(_0886_),
    .Q(\gen_left[0][15] ));
 sky130_fd_sc_hd__dfrtp_2 _4988_ (.CLK(clk),
    .D(_0200_),
    .RESET_B(_0887_),
    .Q(\gen_left[0][16] ));
 sky130_fd_sc_hd__dfrtp_2 _4989_ (.CLK(clk),
    .D(_0201_),
    .RESET_B(_0888_),
    .Q(\gen_left[0][17] ));
 sky130_fd_sc_hd__dfrtp_2 _4990_ (.CLK(clk),
    .D(_0202_),
    .RESET_B(_0889_),
    .Q(\gen_left[0][18] ));
 sky130_fd_sc_hd__dfrtp_2 _4991_ (.CLK(clk),
    .D(_0203_),
    .RESET_B(_0890_),
    .Q(\gen_left[0][19] ));
 sky130_fd_sc_hd__dfrtp_2 _4992_ (.CLK(clk),
    .D(_0205_),
    .RESET_B(_0891_),
    .Q(\gen_left[0][20] ));
 sky130_fd_sc_hd__dfrtp_2 _4993_ (.CLK(clk),
    .D(_0206_),
    .RESET_B(_0892_),
    .Q(\gen_left[0][21] ));
 sky130_fd_sc_hd__dfrtp_2 _4994_ (.CLK(clk),
    .D(_0207_),
    .RESET_B(_0893_),
    .Q(\gen_left[0][22] ));
 sky130_fd_sc_hd__dfrtp_2 _4995_ (.CLK(clk),
    .D(_0208_),
    .RESET_B(_0894_),
    .Q(\gen_left[0][23] ));
 sky130_fd_sc_hd__dfrtp_2 _4996_ (.CLK(clk),
    .D(_0209_),
    .RESET_B(_0895_),
    .Q(\gen_left[0][24] ));
 sky130_fd_sc_hd__dfrtp_2 _4997_ (.CLK(clk),
    .D(_0210_),
    .RESET_B(_0896_),
    .Q(\gen_left[0][25] ));
 sky130_fd_sc_hd__dfrtp_2 _4998_ (.CLK(clk),
    .D(_0211_),
    .RESET_B(_0897_),
    .Q(\gen_left[0][26] ));
 sky130_fd_sc_hd__dfrtp_2 _4999_ (.CLK(clk),
    .D(_0212_),
    .RESET_B(_0898_),
    .Q(\gen_left[0][27] ));
 sky130_fd_sc_hd__dfrtp_2 _5000_ (.CLK(clk),
    .D(_0213_),
    .RESET_B(_0899_),
    .Q(\gen_left[0][28] ));
 sky130_fd_sc_hd__dfrtp_2 _5001_ (.CLK(clk),
    .D(_0214_),
    .RESET_B(_0900_),
    .Q(\gen_left[0][29] ));
 sky130_fd_sc_hd__dfrtp_2 _5002_ (.CLK(clk),
    .D(_0216_),
    .RESET_B(_0901_),
    .Q(\gen_left[0][30] ));
 sky130_fd_sc_hd__dfrtp_2 _5003_ (.CLK(clk),
    .D(_0217_),
    .RESET_B(_0902_),
    .Q(\gen_left[0][31] ));
 sky130_fd_sc_hd__dfrtp_2 _5004_ (.CLK(clk),
    .D(_0321_),
    .RESET_B(_0903_),
    .Q(\gen_left[2][0] ));
 sky130_fd_sc_hd__dfrtp_2 _5005_ (.CLK(clk),
    .D(_0332_),
    .RESET_B(_0904_),
    .Q(\gen_left[2][1] ));
 sky130_fd_sc_hd__dfrtp_2 _5006_ (.CLK(clk),
    .D(_0343_),
    .RESET_B(_0905_),
    .Q(\gen_left[2][2] ));
 sky130_fd_sc_hd__dfrtp_2 _5007_ (.CLK(clk),
    .D(_0346_),
    .RESET_B(_0906_),
    .Q(\gen_left[2][3] ));
 sky130_fd_sc_hd__dfrtp_2 _5008_ (.CLK(clk),
    .D(_0347_),
    .RESET_B(_0907_),
    .Q(\gen_left[2][4] ));
 sky130_fd_sc_hd__dfrtp_2 _5009_ (.CLK(clk),
    .D(_0348_),
    .RESET_B(_0908_),
    .Q(\gen_left[2][5] ));
 sky130_fd_sc_hd__dfrtp_2 _5010_ (.CLK(clk),
    .D(_0349_),
    .RESET_B(_0909_),
    .Q(\gen_left[2][6] ));
 sky130_fd_sc_hd__dfrtp_2 _5011_ (.CLK(clk),
    .D(_0350_),
    .RESET_B(_0910_),
    .Q(\gen_left[2][7] ));
 sky130_fd_sc_hd__dfrtp_2 _5012_ (.CLK(clk),
    .D(_0351_),
    .RESET_B(_0911_),
    .Q(\gen_left[2][8] ));
 sky130_fd_sc_hd__dfrtp_2 _5013_ (.CLK(clk),
    .D(_0352_),
    .RESET_B(_0912_),
    .Q(\gen_left[2][9] ));
 sky130_fd_sc_hd__dfrtp_2 _5014_ (.CLK(clk),
    .D(_0322_),
    .RESET_B(_0913_),
    .Q(\gen_left[2][10] ));
 sky130_fd_sc_hd__dfrtp_2 _5015_ (.CLK(clk),
    .D(_0323_),
    .RESET_B(_0914_),
    .Q(\gen_left[2][11] ));
 sky130_fd_sc_hd__dfrtp_2 _5016_ (.CLK(clk),
    .D(_0324_),
    .RESET_B(_0915_),
    .Q(\gen_left[2][12] ));
 sky130_fd_sc_hd__dfrtp_2 _5017_ (.CLK(clk),
    .D(_0325_),
    .RESET_B(_0916_),
    .Q(\gen_left[2][13] ));
 sky130_fd_sc_hd__dfrtp_2 _5018_ (.CLK(clk),
    .D(_0326_),
    .RESET_B(_0917_),
    .Q(\gen_left[2][14] ));
 sky130_fd_sc_hd__dfrtp_2 _5019_ (.CLK(clk),
    .D(_0327_),
    .RESET_B(_0918_),
    .Q(\gen_left[2][15] ));
 sky130_fd_sc_hd__dfrtp_2 _5020_ (.CLK(clk),
    .D(_0328_),
    .RESET_B(_0919_),
    .Q(\gen_left[2][16] ));
 sky130_fd_sc_hd__dfrtp_2 _5021_ (.CLK(clk),
    .D(_0329_),
    .RESET_B(_0920_),
    .Q(\gen_left[2][17] ));
 sky130_fd_sc_hd__dfrtp_2 _5022_ (.CLK(clk),
    .D(_0330_),
    .RESET_B(_0921_),
    .Q(\gen_left[2][18] ));
 sky130_fd_sc_hd__dfrtp_2 _5023_ (.CLK(clk),
    .D(_0331_),
    .RESET_B(_0922_),
    .Q(\gen_left[2][19] ));
 sky130_fd_sc_hd__dfrtp_2 _5024_ (.CLK(clk),
    .D(_0333_),
    .RESET_B(_0923_),
    .Q(\gen_left[2][20] ));
 sky130_fd_sc_hd__dfrtp_2 _5025_ (.CLK(clk),
    .D(_0334_),
    .RESET_B(_0924_),
    .Q(\gen_left[2][21] ));
 sky130_fd_sc_hd__dfrtp_2 _5026_ (.CLK(clk),
    .D(_0335_),
    .RESET_B(_0925_),
    .Q(\gen_left[2][22] ));
 sky130_fd_sc_hd__dfrtp_2 _5027_ (.CLK(clk),
    .D(_0336_),
    .RESET_B(_0926_),
    .Q(\gen_left[2][23] ));
 sky130_fd_sc_hd__dfrtp_2 _5028_ (.CLK(clk),
    .D(_0337_),
    .RESET_B(_0927_),
    .Q(\gen_left[2][24] ));
 sky130_fd_sc_hd__dfrtp_2 _5029_ (.CLK(clk),
    .D(_0338_),
    .RESET_B(_0928_),
    .Q(\gen_left[2][25] ));
 sky130_fd_sc_hd__dfrtp_2 _5030_ (.CLK(clk),
    .D(_0339_),
    .RESET_B(_0929_),
    .Q(\gen_left[2][26] ));
 sky130_fd_sc_hd__dfrtp_2 _5031_ (.CLK(clk),
    .D(_0340_),
    .RESET_B(_0930_),
    .Q(\gen_left[2][27] ));
 sky130_fd_sc_hd__dfrtp_2 _5032_ (.CLK(clk),
    .D(_0341_),
    .RESET_B(_0931_),
    .Q(\gen_left[2][28] ));
 sky130_fd_sc_hd__dfrtp_2 _5033_ (.CLK(clk),
    .D(_0342_),
    .RESET_B(_0932_),
    .Q(\gen_left[2][29] ));
 sky130_fd_sc_hd__dfrtp_2 _5034_ (.CLK(clk),
    .D(_0344_),
    .RESET_B(_0933_),
    .Q(\gen_left[2][30] ));
 sky130_fd_sc_hd__dfrtp_2 _5035_ (.CLK(clk),
    .D(_0345_),
    .RESET_B(_0934_),
    .Q(\gen_left[2][31] ));
 sky130_fd_sc_hd__dfrtp_2 _5036_ (.CLK(clk),
    .D(_0353_),
    .RESET_B(_0935_),
    .Q(\gen_pe[2].pe_inst.out_right[0] ));
 sky130_fd_sc_hd__dfrtp_2 _5037_ (.CLK(clk),
    .D(_0364_),
    .RESET_B(_0936_),
    .Q(\gen_pe[2].pe_inst.out_right[1] ));
 sky130_fd_sc_hd__dfrtp_2 _5038_ (.CLK(clk),
    .D(_0375_),
    .RESET_B(_0937_),
    .Q(\gen_pe[2].pe_inst.out_right[2] ));
 sky130_fd_sc_hd__dfrtp_2 _5039_ (.CLK(clk),
    .D(_0378_),
    .RESET_B(_0938_),
    .Q(\gen_pe[2].pe_inst.out_right[3] ));
 sky130_fd_sc_hd__dfrtp_2 _5040_ (.CLK(clk),
    .D(_0379_),
    .RESET_B(_0939_),
    .Q(\gen_pe[2].pe_inst.out_right[4] ));
 sky130_fd_sc_hd__dfrtp_2 _5041_ (.CLK(clk),
    .D(_0380_),
    .RESET_B(_0940_),
    .Q(\gen_pe[2].pe_inst.out_right[5] ));
 sky130_fd_sc_hd__dfrtp_2 _5042_ (.CLK(clk),
    .D(_0381_),
    .RESET_B(_0941_),
    .Q(\gen_pe[2].pe_inst.out_right[6] ));
 sky130_fd_sc_hd__dfrtp_2 _5043_ (.CLK(clk),
    .D(_0382_),
    .RESET_B(_0942_),
    .Q(\gen_pe[2].pe_inst.out_right[7] ));
 sky130_fd_sc_hd__dfrtp_2 _5044_ (.CLK(clk),
    .D(_0383_),
    .RESET_B(_0943_),
    .Q(\gen_pe[2].pe_inst.out_right[8] ));
 sky130_fd_sc_hd__dfrtp_2 _5045_ (.CLK(clk),
    .D(_0384_),
    .RESET_B(_0944_),
    .Q(\gen_pe[2].pe_inst.out_right[9] ));
 sky130_fd_sc_hd__dfrtp_2 _5046_ (.CLK(clk),
    .D(_0354_),
    .RESET_B(_0945_),
    .Q(\gen_pe[2].pe_inst.out_right[10] ));
 sky130_fd_sc_hd__dfrtp_2 _5047_ (.CLK(clk),
    .D(_0355_),
    .RESET_B(_0946_),
    .Q(\gen_pe[2].pe_inst.out_right[11] ));
 sky130_fd_sc_hd__dfrtp_2 _5048_ (.CLK(clk),
    .D(_0356_),
    .RESET_B(_0947_),
    .Q(\gen_pe[2].pe_inst.out_right[12] ));
 sky130_fd_sc_hd__dfrtp_2 _5049_ (.CLK(clk),
    .D(_0357_),
    .RESET_B(_0948_),
    .Q(\gen_pe[2].pe_inst.out_right[13] ));
 sky130_fd_sc_hd__dfrtp_2 _5050_ (.CLK(clk),
    .D(_0358_),
    .RESET_B(_0949_),
    .Q(\gen_pe[2].pe_inst.out_right[14] ));
 sky130_fd_sc_hd__dfrtp_2 _5051_ (.CLK(clk),
    .D(_0359_),
    .RESET_B(_0950_),
    .Q(\gen_pe[2].pe_inst.out_right[15] ));
 sky130_fd_sc_hd__dfrtp_2 _5052_ (.CLK(clk),
    .D(_0360_),
    .RESET_B(_0951_),
    .Q(\gen_pe[2].pe_inst.out_right[16] ));
 sky130_fd_sc_hd__dfrtp_2 _5053_ (.CLK(clk),
    .D(_0361_),
    .RESET_B(_0952_),
    .Q(\gen_pe[2].pe_inst.out_right[17] ));
 sky130_fd_sc_hd__dfrtp_2 _5054_ (.CLK(clk),
    .D(_0362_),
    .RESET_B(_0953_),
    .Q(\gen_pe[2].pe_inst.out_right[18] ));
 sky130_fd_sc_hd__dfrtp_2 _5055_ (.CLK(clk),
    .D(_0363_),
    .RESET_B(_0954_),
    .Q(\gen_pe[2].pe_inst.out_right[19] ));
 sky130_fd_sc_hd__dfrtp_2 _5056_ (.CLK(clk),
    .D(_0365_),
    .RESET_B(_0955_),
    .Q(\gen_pe[2].pe_inst.out_right[20] ));
 sky130_fd_sc_hd__dfrtp_2 _5057_ (.CLK(clk),
    .D(_0366_),
    .RESET_B(_0956_),
    .Q(\gen_pe[2].pe_inst.out_right[21] ));
 sky130_fd_sc_hd__dfrtp_2 _5058_ (.CLK(clk),
    .D(_0367_),
    .RESET_B(_0957_),
    .Q(\gen_pe[2].pe_inst.out_right[22] ));
 sky130_fd_sc_hd__dfrtp_2 _5059_ (.CLK(clk),
    .D(_0368_),
    .RESET_B(_0958_),
    .Q(\gen_pe[2].pe_inst.out_right[23] ));
 sky130_fd_sc_hd__dfrtp_2 _5060_ (.CLK(clk),
    .D(_0369_),
    .RESET_B(_0959_),
    .Q(\gen_pe[2].pe_inst.out_right[24] ));
 sky130_fd_sc_hd__dfrtp_2 _5061_ (.CLK(clk),
    .D(_0370_),
    .RESET_B(_0960_),
    .Q(\gen_pe[2].pe_inst.out_right[25] ));
 sky130_fd_sc_hd__dfrtp_2 _5062_ (.CLK(clk),
    .D(_0371_),
    .RESET_B(_0961_),
    .Q(\gen_pe[2].pe_inst.out_right[26] ));
 sky130_fd_sc_hd__dfrtp_2 _5063_ (.CLK(clk),
    .D(_0372_),
    .RESET_B(_0962_),
    .Q(\gen_pe[2].pe_inst.out_right[27] ));
 sky130_fd_sc_hd__dfrtp_2 _5064_ (.CLK(clk),
    .D(_0373_),
    .RESET_B(_0963_),
    .Q(\gen_pe[2].pe_inst.out_right[28] ));
 sky130_fd_sc_hd__dfrtp_2 _5065_ (.CLK(clk),
    .D(_0374_),
    .RESET_B(_0964_),
    .Q(\gen_pe[2].pe_inst.out_right[29] ));
 sky130_fd_sc_hd__dfrtp_2 _5066_ (.CLK(clk),
    .D(_0376_),
    .RESET_B(_0965_),
    .Q(\gen_pe[2].pe_inst.out_right[30] ));
 sky130_fd_sc_hd__dfrtp_2 _5067_ (.CLK(clk),
    .D(_0377_),
    .RESET_B(_0966_),
    .Q(\gen_pe[2].pe_inst.out_right[31] ));
 sky130_fd_sc_hd__dfrtp_2 _5068_ (.CLK(clk),
    .D(_0513_),
    .RESET_B(_0967_),
    .Q(\gen_left[5][0] ));
 sky130_fd_sc_hd__dfrtp_2 _5069_ (.CLK(clk),
    .D(_0524_),
    .RESET_B(_0968_),
    .Q(\gen_left[5][1] ));
 sky130_fd_sc_hd__dfrtp_2 _5070_ (.CLK(clk),
    .D(_0535_),
    .RESET_B(_0969_),
    .Q(\gen_left[5][2] ));
 sky130_fd_sc_hd__dfrtp_2 _5071_ (.CLK(clk),
    .D(_0538_),
    .RESET_B(_0970_),
    .Q(\gen_left[5][3] ));
 sky130_fd_sc_hd__dfrtp_2 _5072_ (.CLK(clk),
    .D(_0539_),
    .RESET_B(_0971_),
    .Q(\gen_left[5][4] ));
 sky130_fd_sc_hd__dfrtp_2 _5073_ (.CLK(clk),
    .D(_0540_),
    .RESET_B(_0972_),
    .Q(\gen_left[5][5] ));
 sky130_fd_sc_hd__dfrtp_2 _5074_ (.CLK(clk),
    .D(_0541_),
    .RESET_B(_0973_),
    .Q(\gen_left[5][6] ));
 sky130_fd_sc_hd__dfrtp_2 _5075_ (.CLK(clk),
    .D(_0542_),
    .RESET_B(_0974_),
    .Q(\gen_left[5][7] ));
 sky130_fd_sc_hd__dfrtp_2 _5076_ (.CLK(clk),
    .D(_0543_),
    .RESET_B(_0975_),
    .Q(\gen_left[5][8] ));
 sky130_fd_sc_hd__dfrtp_2 _5077_ (.CLK(clk),
    .D(_0544_),
    .RESET_B(_0976_),
    .Q(\gen_left[5][9] ));
 sky130_fd_sc_hd__dfrtp_2 _5078_ (.CLK(clk),
    .D(_0514_),
    .RESET_B(_0977_),
    .Q(\gen_left[5][10] ));
 sky130_fd_sc_hd__dfrtp_2 _5079_ (.CLK(clk),
    .D(_0515_),
    .RESET_B(_0978_),
    .Q(\gen_left[5][11] ));
 sky130_fd_sc_hd__dfrtp_2 _5080_ (.CLK(clk),
    .D(_0516_),
    .RESET_B(_0979_),
    .Q(\gen_left[5][12] ));
 sky130_fd_sc_hd__dfrtp_2 _5081_ (.CLK(clk),
    .D(_0517_),
    .RESET_B(_0980_),
    .Q(\gen_left[5][13] ));
 sky130_fd_sc_hd__dfrtp_2 _5082_ (.CLK(clk),
    .D(_0518_),
    .RESET_B(_0981_),
    .Q(\gen_left[5][14] ));
 sky130_fd_sc_hd__dfrtp_2 _5083_ (.CLK(clk),
    .D(_0519_),
    .RESET_B(_0982_),
    .Q(\gen_left[5][15] ));
 sky130_fd_sc_hd__dfrtp_2 _5084_ (.CLK(clk),
    .D(_0520_),
    .RESET_B(_0983_),
    .Q(\gen_left[5][16] ));
 sky130_fd_sc_hd__dfrtp_2 _5085_ (.CLK(clk),
    .D(_0521_),
    .RESET_B(_0984_),
    .Q(\gen_left[5][17] ));
 sky130_fd_sc_hd__dfrtp_2 _5086_ (.CLK(clk),
    .D(_0522_),
    .RESET_B(_0985_),
    .Q(\gen_left[5][18] ));
 sky130_fd_sc_hd__dfrtp_2 _5087_ (.CLK(clk),
    .D(_0523_),
    .RESET_B(_0986_),
    .Q(\gen_left[5][19] ));
 sky130_fd_sc_hd__dfrtp_2 _5088_ (.CLK(clk),
    .D(_0525_),
    .RESET_B(_0987_),
    .Q(\gen_left[5][20] ));
 sky130_fd_sc_hd__dfrtp_2 _5089_ (.CLK(clk),
    .D(_0526_),
    .RESET_B(_0988_),
    .Q(\gen_left[5][21] ));
 sky130_fd_sc_hd__dfrtp_2 _5090_ (.CLK(clk),
    .D(_0527_),
    .RESET_B(_0989_),
    .Q(\gen_left[5][22] ));
 sky130_fd_sc_hd__dfrtp_2 _5091_ (.CLK(clk),
    .D(_0528_),
    .RESET_B(_0990_),
    .Q(\gen_left[5][23] ));
 sky130_fd_sc_hd__dfrtp_2 _5092_ (.CLK(clk),
    .D(_0529_),
    .RESET_B(_0991_),
    .Q(\gen_left[5][24] ));
 sky130_fd_sc_hd__dfrtp_2 _5093_ (.CLK(clk),
    .D(_0530_),
    .RESET_B(_0992_),
    .Q(\gen_left[5][25] ));
 sky130_fd_sc_hd__dfrtp_2 _5094_ (.CLK(clk),
    .D(_0531_),
    .RESET_B(_0993_),
    .Q(\gen_left[5][26] ));
 sky130_fd_sc_hd__dfrtp_2 _5095_ (.CLK(clk),
    .D(_0532_),
    .RESET_B(_0994_),
    .Q(\gen_left[5][27] ));
 sky130_fd_sc_hd__dfrtp_2 _5096_ (.CLK(clk),
    .D(_0533_),
    .RESET_B(_0995_),
    .Q(\gen_left[5][28] ));
 sky130_fd_sc_hd__dfrtp_2 _5097_ (.CLK(clk),
    .D(_0534_),
    .RESET_B(_0996_),
    .Q(\gen_left[5][29] ));
 sky130_fd_sc_hd__dfrtp_2 _5098_ (.CLK(clk),
    .D(_0536_),
    .RESET_B(_0997_),
    .Q(\gen_left[5][30] ));
 sky130_fd_sc_hd__dfrtp_2 _5099_ (.CLK(clk),
    .D(_0537_),
    .RESET_B(_0998_),
    .Q(\gen_left[5][31] ));
 sky130_fd_sc_hd__dfrtp_2 _5100_ (.CLK(clk),
    .D(_0545_),
    .RESET_B(_0999_),
    .Q(\gen_pe[5].pe_inst.out_right[0] ));
 sky130_fd_sc_hd__dfrtp_2 _5101_ (.CLK(clk),
    .D(_0556_),
    .RESET_B(_1000_),
    .Q(\gen_pe[5].pe_inst.out_right[1] ));
 sky130_fd_sc_hd__dfrtp_2 _5102_ (.CLK(clk),
    .D(_0567_),
    .RESET_B(_1001_),
    .Q(\gen_pe[5].pe_inst.out_right[2] ));
 sky130_fd_sc_hd__dfrtp_2 _5103_ (.CLK(clk),
    .D(_0570_),
    .RESET_B(_1002_),
    .Q(\gen_pe[5].pe_inst.out_right[3] ));
 sky130_fd_sc_hd__dfrtp_2 _5104_ (.CLK(clk),
    .D(_0571_),
    .RESET_B(_1003_),
    .Q(\gen_pe[5].pe_inst.out_right[4] ));
 sky130_fd_sc_hd__dfrtp_2 _5105_ (.CLK(clk),
    .D(_0572_),
    .RESET_B(_1004_),
    .Q(\gen_pe[5].pe_inst.out_right[5] ));
 sky130_fd_sc_hd__dfrtp_2 _5106_ (.CLK(clk),
    .D(_0573_),
    .RESET_B(_1005_),
    .Q(\gen_pe[5].pe_inst.out_right[6] ));
 sky130_fd_sc_hd__dfrtp_2 _5107_ (.CLK(clk),
    .D(_0574_),
    .RESET_B(_1006_),
    .Q(\gen_pe[5].pe_inst.out_right[7] ));
 sky130_fd_sc_hd__dfrtp_2 _5108_ (.CLK(clk),
    .D(_0575_),
    .RESET_B(_1007_),
    .Q(\gen_pe[5].pe_inst.out_right[8] ));
 sky130_fd_sc_hd__dfrtp_2 _5109_ (.CLK(clk),
    .D(_0576_),
    .RESET_B(_1008_),
    .Q(\gen_pe[5].pe_inst.out_right[9] ));
 sky130_fd_sc_hd__dfrtp_2 _5110_ (.CLK(clk),
    .D(_0546_),
    .RESET_B(_1009_),
    .Q(\gen_pe[5].pe_inst.out_right[10] ));
 sky130_fd_sc_hd__dfrtp_2 _5111_ (.CLK(clk),
    .D(_0547_),
    .RESET_B(_1010_),
    .Q(\gen_pe[5].pe_inst.out_right[11] ));
 sky130_fd_sc_hd__dfrtp_2 _5112_ (.CLK(clk),
    .D(_0548_),
    .RESET_B(_1011_),
    .Q(\gen_pe[5].pe_inst.out_right[12] ));
 sky130_fd_sc_hd__dfrtp_2 _5113_ (.CLK(clk),
    .D(_0549_),
    .RESET_B(_1012_),
    .Q(\gen_pe[5].pe_inst.out_right[13] ));
 sky130_fd_sc_hd__dfrtp_2 _5114_ (.CLK(clk),
    .D(_0550_),
    .RESET_B(_1013_),
    .Q(\gen_pe[5].pe_inst.out_right[14] ));
 sky130_fd_sc_hd__dfrtp_2 _5115_ (.CLK(clk),
    .D(_0551_),
    .RESET_B(_1014_),
    .Q(\gen_pe[5].pe_inst.out_right[15] ));
 sky130_fd_sc_hd__dfrtp_2 _5116_ (.CLK(clk),
    .D(_0552_),
    .RESET_B(_1015_),
    .Q(\gen_pe[5].pe_inst.out_right[16] ));
 sky130_fd_sc_hd__dfrtp_2 _5117_ (.CLK(clk),
    .D(_0553_),
    .RESET_B(_1016_),
    .Q(\gen_pe[5].pe_inst.out_right[17] ));
 sky130_fd_sc_hd__dfrtp_2 _5118_ (.CLK(clk),
    .D(_0554_),
    .RESET_B(_1017_),
    .Q(\gen_pe[5].pe_inst.out_right[18] ));
 sky130_fd_sc_hd__dfrtp_2 _5119_ (.CLK(clk),
    .D(_0555_),
    .RESET_B(_1018_),
    .Q(\gen_pe[5].pe_inst.out_right[19] ));
 sky130_fd_sc_hd__dfrtp_2 _5120_ (.CLK(clk),
    .D(_0557_),
    .RESET_B(_1019_),
    .Q(\gen_pe[5].pe_inst.out_right[20] ));
 sky130_fd_sc_hd__dfrtp_2 _5121_ (.CLK(clk),
    .D(_0558_),
    .RESET_B(_1020_),
    .Q(\gen_pe[5].pe_inst.out_right[21] ));
 sky130_fd_sc_hd__dfrtp_2 _5122_ (.CLK(clk),
    .D(_0559_),
    .RESET_B(_1021_),
    .Q(\gen_pe[5].pe_inst.out_right[22] ));
 sky130_fd_sc_hd__dfrtp_2 _5123_ (.CLK(clk),
    .D(_0560_),
    .RESET_B(_1022_),
    .Q(\gen_pe[5].pe_inst.out_right[23] ));
 sky130_fd_sc_hd__dfrtp_2 _5124_ (.CLK(clk),
    .D(_0561_),
    .RESET_B(_1023_),
    .Q(\gen_pe[5].pe_inst.out_right[24] ));
 sky130_fd_sc_hd__dfrtp_2 _5125_ (.CLK(clk),
    .D(_0562_),
    .RESET_B(_1024_),
    .Q(\gen_pe[5].pe_inst.out_right[25] ));
 sky130_fd_sc_hd__dfrtp_2 _5126_ (.CLK(clk),
    .D(_0563_),
    .RESET_B(_1025_),
    .Q(\gen_pe[5].pe_inst.out_right[26] ));
 sky130_fd_sc_hd__dfrtp_2 _5127_ (.CLK(clk),
    .D(_0564_),
    .RESET_B(_1026_),
    .Q(\gen_pe[5].pe_inst.out_right[27] ));
 sky130_fd_sc_hd__dfrtp_2 _5128_ (.CLK(clk),
    .D(_0565_),
    .RESET_B(_1027_),
    .Q(\gen_pe[5].pe_inst.out_right[28] ));
 sky130_fd_sc_hd__dfrtp_2 _5129_ (.CLK(clk),
    .D(_0566_),
    .RESET_B(_1028_),
    .Q(\gen_pe[5].pe_inst.out_right[29] ));
 sky130_fd_sc_hd__dfrtp_2 _5130_ (.CLK(clk),
    .D(_0568_),
    .RESET_B(_1029_),
    .Q(\gen_pe[5].pe_inst.out_right[30] ));
 sky130_fd_sc_hd__dfrtp_2 _5131_ (.CLK(clk),
    .D(_0569_),
    .RESET_B(_1030_),
    .Q(\gen_pe[5].pe_inst.out_right[31] ));
 sky130_fd_sc_hd__dfrtp_2 _5132_ (.CLK(clk),
    .D(_0449_),
    .RESET_B(_1031_),
    .Q(\gen_left[4][0] ));
 sky130_fd_sc_hd__dfrtp_2 _5133_ (.CLK(clk),
    .D(_0460_),
    .RESET_B(_1032_),
    .Q(\gen_left[4][1] ));
 sky130_fd_sc_hd__dfrtp_2 _5134_ (.CLK(clk),
    .D(_0471_),
    .RESET_B(_1033_),
    .Q(\gen_left[4][2] ));
 sky130_fd_sc_hd__dfrtp_2 _5135_ (.CLK(clk),
    .D(_0474_),
    .RESET_B(_1034_),
    .Q(\gen_left[4][3] ));
 sky130_fd_sc_hd__dfrtp_2 _5136_ (.CLK(clk),
    .D(_0475_),
    .RESET_B(_1035_),
    .Q(\gen_left[4][4] ));
 sky130_fd_sc_hd__dfrtp_2 _5137_ (.CLK(clk),
    .D(_0476_),
    .RESET_B(_1036_),
    .Q(\gen_left[4][5] ));
 sky130_fd_sc_hd__dfrtp_2 _5138_ (.CLK(clk),
    .D(_0477_),
    .RESET_B(_1037_),
    .Q(\gen_left[4][6] ));
 sky130_fd_sc_hd__dfrtp_2 _5139_ (.CLK(clk),
    .D(_0478_),
    .RESET_B(_1038_),
    .Q(\gen_left[4][7] ));
 sky130_fd_sc_hd__dfrtp_2 _5140_ (.CLK(clk),
    .D(_0479_),
    .RESET_B(_1039_),
    .Q(\gen_left[4][8] ));
 sky130_fd_sc_hd__dfrtp_2 _5141_ (.CLK(clk),
    .D(_0480_),
    .RESET_B(_1040_),
    .Q(\gen_left[4][9] ));
 sky130_fd_sc_hd__dfrtp_2 _5142_ (.CLK(clk),
    .D(_0450_),
    .RESET_B(_1041_),
    .Q(\gen_left[4][10] ));
 sky130_fd_sc_hd__dfrtp_2 _5143_ (.CLK(clk),
    .D(_0451_),
    .RESET_B(_1042_),
    .Q(\gen_left[4][11] ));
 sky130_fd_sc_hd__dfrtp_2 _5144_ (.CLK(clk),
    .D(_0452_),
    .RESET_B(_1043_),
    .Q(\gen_left[4][12] ));
 sky130_fd_sc_hd__dfrtp_2 _5145_ (.CLK(clk),
    .D(_0453_),
    .RESET_B(_1044_),
    .Q(\gen_left[4][13] ));
 sky130_fd_sc_hd__dfrtp_2 _5146_ (.CLK(clk),
    .D(_0454_),
    .RESET_B(_1045_),
    .Q(\gen_left[4][14] ));
 sky130_fd_sc_hd__dfrtp_2 _5147_ (.CLK(clk),
    .D(_0455_),
    .RESET_B(_1046_),
    .Q(\gen_left[4][15] ));
 sky130_fd_sc_hd__dfrtp_2 _5148_ (.CLK(clk),
    .D(_0456_),
    .RESET_B(_1047_),
    .Q(\gen_left[4][16] ));
 sky130_fd_sc_hd__dfrtp_2 _5149_ (.CLK(clk),
    .D(_0457_),
    .RESET_B(_1048_),
    .Q(\gen_left[4][17] ));
 sky130_fd_sc_hd__dfrtp_2 _5150_ (.CLK(clk),
    .D(_0458_),
    .RESET_B(_1049_),
    .Q(\gen_left[4][18] ));
 sky130_fd_sc_hd__dfrtp_2 _5151_ (.CLK(clk),
    .D(_0459_),
    .RESET_B(_1050_),
    .Q(\gen_left[4][19] ));
 sky130_fd_sc_hd__dfrtp_2 _5152_ (.CLK(clk),
    .D(_0461_),
    .RESET_B(_1051_),
    .Q(\gen_left[4][20] ));
 sky130_fd_sc_hd__dfrtp_2 _5153_ (.CLK(clk),
    .D(_0462_),
    .RESET_B(_1052_),
    .Q(\gen_left[4][21] ));
 sky130_fd_sc_hd__dfrtp_2 _5154_ (.CLK(clk),
    .D(_0463_),
    .RESET_B(_1053_),
    .Q(\gen_left[4][22] ));
 sky130_fd_sc_hd__dfrtp_2 _5155_ (.CLK(clk),
    .D(_0464_),
    .RESET_B(_1054_),
    .Q(\gen_left[4][23] ));
 sky130_fd_sc_hd__dfrtp_2 _5156_ (.CLK(clk),
    .D(_0465_),
    .RESET_B(_1055_),
    .Q(\gen_left[4][24] ));
 sky130_fd_sc_hd__dfrtp_2 _5157_ (.CLK(clk),
    .D(_0466_),
    .RESET_B(_1056_),
    .Q(\gen_left[4][25] ));
 sky130_fd_sc_hd__dfrtp_2 _5158_ (.CLK(clk),
    .D(_0467_),
    .RESET_B(_1057_),
    .Q(\gen_left[4][26] ));
 sky130_fd_sc_hd__dfrtp_2 _5159_ (.CLK(clk),
    .D(_0468_),
    .RESET_B(_1058_),
    .Q(\gen_left[4][27] ));
 sky130_fd_sc_hd__dfrtp_2 _5160_ (.CLK(clk),
    .D(_0469_),
    .RESET_B(_1059_),
    .Q(\gen_left[4][28] ));
 sky130_fd_sc_hd__dfrtp_2 _5161_ (.CLK(clk),
    .D(_0470_),
    .RESET_B(_1060_),
    .Q(\gen_left[4][29] ));
 sky130_fd_sc_hd__dfrtp_2 _5162_ (.CLK(clk),
    .D(_0472_),
    .RESET_B(_1061_),
    .Q(\gen_left[4][30] ));
 sky130_fd_sc_hd__dfrtp_2 _5163_ (.CLK(clk),
    .D(_0473_),
    .RESET_B(_1062_),
    .Q(\gen_left[4][31] ));
 sky130_fd_sc_hd__dfrtp_2 _5164_ (.CLK(clk),
    .D(_0481_),
    .RESET_B(_1063_),
    .Q(\gen_pe[4].pe_inst.out_right[0] ));
 sky130_fd_sc_hd__dfrtp_2 _5165_ (.CLK(clk),
    .D(_0492_),
    .RESET_B(_1064_),
    .Q(\gen_pe[4].pe_inst.out_right[1] ));
 sky130_fd_sc_hd__dfrtp_2 _5166_ (.CLK(clk),
    .D(_0503_),
    .RESET_B(_1065_),
    .Q(\gen_pe[4].pe_inst.out_right[2] ));
 sky130_fd_sc_hd__dfrtp_2 _5167_ (.CLK(clk),
    .D(_0506_),
    .RESET_B(_1066_),
    .Q(\gen_pe[4].pe_inst.out_right[3] ));
 sky130_fd_sc_hd__dfrtp_2 _5168_ (.CLK(clk),
    .D(_0507_),
    .RESET_B(_1067_),
    .Q(\gen_pe[4].pe_inst.out_right[4] ));
 sky130_fd_sc_hd__dfrtp_2 _5169_ (.CLK(clk),
    .D(_0508_),
    .RESET_B(_1068_),
    .Q(\gen_pe[4].pe_inst.out_right[5] ));
 sky130_fd_sc_hd__dfrtp_2 _5170_ (.CLK(clk),
    .D(_0509_),
    .RESET_B(_1069_),
    .Q(\gen_pe[4].pe_inst.out_right[6] ));
 sky130_fd_sc_hd__dfrtp_2 _5171_ (.CLK(clk),
    .D(_0510_),
    .RESET_B(_1070_),
    .Q(\gen_pe[4].pe_inst.out_right[7] ));
 sky130_fd_sc_hd__dfrtp_2 _5172_ (.CLK(clk),
    .D(_0511_),
    .RESET_B(_1071_),
    .Q(\gen_pe[4].pe_inst.out_right[8] ));
 sky130_fd_sc_hd__dfrtp_2 _5173_ (.CLK(clk),
    .D(_0512_),
    .RESET_B(_1072_),
    .Q(\gen_pe[4].pe_inst.out_right[9] ));
 sky130_fd_sc_hd__dfrtp_2 _5174_ (.CLK(clk),
    .D(_0482_),
    .RESET_B(_1073_),
    .Q(\gen_pe[4].pe_inst.out_right[10] ));
 sky130_fd_sc_hd__dfrtp_2 _5175_ (.CLK(clk),
    .D(_0483_),
    .RESET_B(_1074_),
    .Q(\gen_pe[4].pe_inst.out_right[11] ));
 sky130_fd_sc_hd__dfrtp_2 _5176_ (.CLK(clk),
    .D(_0484_),
    .RESET_B(_1075_),
    .Q(\gen_pe[4].pe_inst.out_right[12] ));
 sky130_fd_sc_hd__dfrtp_2 _5177_ (.CLK(clk),
    .D(_0485_),
    .RESET_B(_1076_),
    .Q(\gen_pe[4].pe_inst.out_right[13] ));
 sky130_fd_sc_hd__dfrtp_2 _5178_ (.CLK(clk),
    .D(_0486_),
    .RESET_B(_1077_),
    .Q(\gen_pe[4].pe_inst.out_right[14] ));
 sky130_fd_sc_hd__dfrtp_2 _5179_ (.CLK(clk),
    .D(_0487_),
    .RESET_B(_1078_),
    .Q(\gen_pe[4].pe_inst.out_right[15] ));
 sky130_fd_sc_hd__dfrtp_2 _5180_ (.CLK(clk),
    .D(_0488_),
    .RESET_B(_1079_),
    .Q(\gen_pe[4].pe_inst.out_right[16] ));
 sky130_fd_sc_hd__dfrtp_2 _5181_ (.CLK(clk),
    .D(_0489_),
    .RESET_B(_1080_),
    .Q(\gen_pe[4].pe_inst.out_right[17] ));
 sky130_fd_sc_hd__dfrtp_2 _5182_ (.CLK(clk),
    .D(_0490_),
    .RESET_B(_1081_),
    .Q(\gen_pe[4].pe_inst.out_right[18] ));
 sky130_fd_sc_hd__dfrtp_2 _5183_ (.CLK(clk),
    .D(_0491_),
    .RESET_B(_1082_),
    .Q(\gen_pe[4].pe_inst.out_right[19] ));
 sky130_fd_sc_hd__dfrtp_2 _5184_ (.CLK(clk),
    .D(_0493_),
    .RESET_B(_1083_),
    .Q(\gen_pe[4].pe_inst.out_right[20] ));
 sky130_fd_sc_hd__dfrtp_2 _5185_ (.CLK(clk),
    .D(_0494_),
    .RESET_B(_1084_),
    .Q(\gen_pe[4].pe_inst.out_right[21] ));
 sky130_fd_sc_hd__dfrtp_2 _5186_ (.CLK(clk),
    .D(_0495_),
    .RESET_B(_1085_),
    .Q(\gen_pe[4].pe_inst.out_right[22] ));
 sky130_fd_sc_hd__dfrtp_2 _5187_ (.CLK(clk),
    .D(_0496_),
    .RESET_B(_1086_),
    .Q(\gen_pe[4].pe_inst.out_right[23] ));
 sky130_fd_sc_hd__dfrtp_2 _5188_ (.CLK(clk),
    .D(_0497_),
    .RESET_B(_1087_),
    .Q(\gen_pe[4].pe_inst.out_right[24] ));
 sky130_fd_sc_hd__dfrtp_2 _5189_ (.CLK(clk),
    .D(_0498_),
    .RESET_B(_1088_),
    .Q(\gen_pe[4].pe_inst.out_right[25] ));
 sky130_fd_sc_hd__dfrtp_2 _5190_ (.CLK(clk),
    .D(_0499_),
    .RESET_B(_1089_),
    .Q(\gen_pe[4].pe_inst.out_right[26] ));
 sky130_fd_sc_hd__dfrtp_2 _5191_ (.CLK(clk),
    .D(_0500_),
    .RESET_B(_1090_),
    .Q(\gen_pe[4].pe_inst.out_right[27] ));
 sky130_fd_sc_hd__dfrtp_2 _5192_ (.CLK(clk),
    .D(_0501_),
    .RESET_B(_1091_),
    .Q(\gen_pe[4].pe_inst.out_right[28] ));
 sky130_fd_sc_hd__dfrtp_2 _5193_ (.CLK(clk),
    .D(_0502_),
    .RESET_B(_1092_),
    .Q(\gen_pe[4].pe_inst.out_right[29] ));
 sky130_fd_sc_hd__dfrtp_2 _5194_ (.CLK(clk),
    .D(_0504_),
    .RESET_B(_1093_),
    .Q(\gen_pe[4].pe_inst.out_right[30] ));
 sky130_fd_sc_hd__dfrtp_2 _5195_ (.CLK(clk),
    .D(_0505_),
    .RESET_B(_1094_),
    .Q(\gen_pe[4].pe_inst.out_right[31] ));
 sky130_fd_sc_hd__dfrtp_2 _5196_ (.CLK(clk),
    .D(_0385_),
    .RESET_B(_1095_),
    .Q(\gen_left[3][0] ));
 sky130_fd_sc_hd__dfrtp_2 _5197_ (.CLK(clk),
    .D(_0396_),
    .RESET_B(_1096_),
    .Q(\gen_left[3][1] ));
 sky130_fd_sc_hd__dfrtp_2 _5198_ (.CLK(clk),
    .D(_0407_),
    .RESET_B(_1097_),
    .Q(\gen_left[3][2] ));
 sky130_fd_sc_hd__dfrtp_2 _5199_ (.CLK(clk),
    .D(_0410_),
    .RESET_B(_1098_),
    .Q(\gen_left[3][3] ));
 sky130_fd_sc_hd__dfrtp_2 _5200_ (.CLK(clk),
    .D(_0411_),
    .RESET_B(_1099_),
    .Q(\gen_left[3][4] ));
 sky130_fd_sc_hd__dfrtp_2 _5201_ (.CLK(clk),
    .D(_0412_),
    .RESET_B(_1100_),
    .Q(\gen_left[3][5] ));
 sky130_fd_sc_hd__dfrtp_2 _5202_ (.CLK(clk),
    .D(_0413_),
    .RESET_B(_1101_),
    .Q(\gen_left[3][6] ));
 sky130_fd_sc_hd__dfrtp_2 _5203_ (.CLK(clk),
    .D(_0414_),
    .RESET_B(_1102_),
    .Q(\gen_left[3][7] ));
 sky130_fd_sc_hd__dfrtp_2 _5204_ (.CLK(clk),
    .D(_0415_),
    .RESET_B(_1103_),
    .Q(\gen_left[3][8] ));
 sky130_fd_sc_hd__dfrtp_2 _5205_ (.CLK(clk),
    .D(_0416_),
    .RESET_B(_1104_),
    .Q(\gen_left[3][9] ));
 sky130_fd_sc_hd__dfrtp_2 _5206_ (.CLK(clk),
    .D(_0386_),
    .RESET_B(_1105_),
    .Q(\gen_left[3][10] ));
 sky130_fd_sc_hd__dfrtp_2 _5207_ (.CLK(clk),
    .D(_0387_),
    .RESET_B(_1106_),
    .Q(\gen_left[3][11] ));
 sky130_fd_sc_hd__dfrtp_2 _5208_ (.CLK(clk),
    .D(_0388_),
    .RESET_B(_1107_),
    .Q(\gen_left[3][12] ));
 sky130_fd_sc_hd__dfrtp_2 _5209_ (.CLK(clk),
    .D(_0389_),
    .RESET_B(_1108_),
    .Q(\gen_left[3][13] ));
 sky130_fd_sc_hd__dfrtp_2 _5210_ (.CLK(clk),
    .D(_0390_),
    .RESET_B(_1109_),
    .Q(\gen_left[3][14] ));
 sky130_fd_sc_hd__dfrtp_2 _5211_ (.CLK(clk),
    .D(_0391_),
    .RESET_B(_1110_),
    .Q(\gen_left[3][15] ));
 sky130_fd_sc_hd__dfrtp_2 _5212_ (.CLK(clk),
    .D(_0392_),
    .RESET_B(_1111_),
    .Q(\gen_left[3][16] ));
 sky130_fd_sc_hd__dfrtp_2 _5213_ (.CLK(clk),
    .D(_0393_),
    .RESET_B(_1112_),
    .Q(\gen_left[3][17] ));
 sky130_fd_sc_hd__dfrtp_2 _5214_ (.CLK(clk),
    .D(_0394_),
    .RESET_B(_1113_),
    .Q(\gen_left[3][18] ));
 sky130_fd_sc_hd__dfrtp_2 _5215_ (.CLK(clk),
    .D(_0395_),
    .RESET_B(_1114_),
    .Q(\gen_left[3][19] ));
 sky130_fd_sc_hd__dfrtp_2 _5216_ (.CLK(clk),
    .D(_0397_),
    .RESET_B(_1115_),
    .Q(\gen_left[3][20] ));
 sky130_fd_sc_hd__dfrtp_2 _5217_ (.CLK(clk),
    .D(_0398_),
    .RESET_B(_1116_),
    .Q(\gen_left[3][21] ));
 sky130_fd_sc_hd__dfrtp_2 _5218_ (.CLK(clk),
    .D(_0399_),
    .RESET_B(_1117_),
    .Q(\gen_left[3][22] ));
 sky130_fd_sc_hd__dfrtp_2 _5219_ (.CLK(clk),
    .D(_0400_),
    .RESET_B(_1118_),
    .Q(\gen_left[3][23] ));
 sky130_fd_sc_hd__dfrtp_2 _5220_ (.CLK(clk),
    .D(_0401_),
    .RESET_B(_1119_),
    .Q(\gen_left[3][24] ));
 sky130_fd_sc_hd__dfrtp_2 _5221_ (.CLK(clk),
    .D(_0402_),
    .RESET_B(_1120_),
    .Q(\gen_left[3][25] ));
 sky130_fd_sc_hd__dfrtp_2 _5222_ (.CLK(clk),
    .D(_0403_),
    .RESET_B(_1121_),
    .Q(\gen_left[3][26] ));
 sky130_fd_sc_hd__dfrtp_2 _5223_ (.CLK(clk),
    .D(_0404_),
    .RESET_B(_1122_),
    .Q(\gen_left[3][27] ));
 sky130_fd_sc_hd__dfrtp_2 _5224_ (.CLK(clk),
    .D(_0405_),
    .RESET_B(_1123_),
    .Q(\gen_left[3][28] ));
 sky130_fd_sc_hd__dfrtp_2 _5225_ (.CLK(clk),
    .D(_0406_),
    .RESET_B(_1124_),
    .Q(\gen_left[3][29] ));
 sky130_fd_sc_hd__dfrtp_2 _5226_ (.CLK(clk),
    .D(_0408_),
    .RESET_B(_1125_),
    .Q(\gen_left[3][30] ));
 sky130_fd_sc_hd__dfrtp_2 _5227_ (.CLK(clk),
    .D(_0409_),
    .RESET_B(_1126_),
    .Q(\gen_left[3][31] ));
 sky130_fd_sc_hd__dfrtp_2 _5228_ (.CLK(clk),
    .D(_0417_),
    .RESET_B(_1127_),
    .Q(\gen_pe[3].pe_inst.out_right[0] ));
 sky130_fd_sc_hd__dfrtp_2 _5229_ (.CLK(clk),
    .D(_0428_),
    .RESET_B(_1128_),
    .Q(\gen_pe[3].pe_inst.out_right[1] ));
 sky130_fd_sc_hd__dfrtp_2 _5230_ (.CLK(clk),
    .D(_0439_),
    .RESET_B(_1129_),
    .Q(\gen_pe[3].pe_inst.out_right[2] ));
 sky130_fd_sc_hd__dfrtp_2 _5231_ (.CLK(clk),
    .D(_0442_),
    .RESET_B(_1130_),
    .Q(\gen_pe[3].pe_inst.out_right[3] ));
 sky130_fd_sc_hd__dfrtp_2 _5232_ (.CLK(clk),
    .D(_0443_),
    .RESET_B(_1131_),
    .Q(\gen_pe[3].pe_inst.out_right[4] ));
 sky130_fd_sc_hd__dfrtp_2 _5233_ (.CLK(clk),
    .D(_0444_),
    .RESET_B(_1132_),
    .Q(\gen_pe[3].pe_inst.out_right[5] ));
 sky130_fd_sc_hd__dfrtp_2 _5234_ (.CLK(clk),
    .D(_0445_),
    .RESET_B(_1133_),
    .Q(\gen_pe[3].pe_inst.out_right[6] ));
 sky130_fd_sc_hd__dfrtp_2 _5235_ (.CLK(clk),
    .D(_0446_),
    .RESET_B(_1134_),
    .Q(\gen_pe[3].pe_inst.out_right[7] ));
 sky130_fd_sc_hd__dfrtp_2 _5236_ (.CLK(clk),
    .D(_0447_),
    .RESET_B(_1135_),
    .Q(\gen_pe[3].pe_inst.out_right[8] ));
 sky130_fd_sc_hd__dfrtp_2 _5237_ (.CLK(clk),
    .D(_0448_),
    .RESET_B(_1136_),
    .Q(\gen_pe[3].pe_inst.out_right[9] ));
 sky130_fd_sc_hd__dfrtp_2 _5238_ (.CLK(clk),
    .D(_0418_),
    .RESET_B(_1137_),
    .Q(\gen_pe[3].pe_inst.out_right[10] ));
 sky130_fd_sc_hd__dfrtp_2 _5239_ (.CLK(clk),
    .D(_0419_),
    .RESET_B(_1138_),
    .Q(\gen_pe[3].pe_inst.out_right[11] ));
 sky130_fd_sc_hd__dfrtp_2 _5240_ (.CLK(clk),
    .D(_0420_),
    .RESET_B(_1139_),
    .Q(\gen_pe[3].pe_inst.out_right[12] ));
 sky130_fd_sc_hd__dfrtp_2 _5241_ (.CLK(clk),
    .D(_0421_),
    .RESET_B(_1140_),
    .Q(\gen_pe[3].pe_inst.out_right[13] ));
 sky130_fd_sc_hd__dfrtp_2 _5242_ (.CLK(clk),
    .D(_0422_),
    .RESET_B(_1141_),
    .Q(\gen_pe[3].pe_inst.out_right[14] ));
 sky130_fd_sc_hd__dfrtp_2 _5243_ (.CLK(clk),
    .D(_0423_),
    .RESET_B(_1142_),
    .Q(\gen_pe[3].pe_inst.out_right[15] ));
 sky130_fd_sc_hd__dfrtp_2 _5244_ (.CLK(clk),
    .D(_0424_),
    .RESET_B(_1143_),
    .Q(\gen_pe[3].pe_inst.out_right[16] ));
 sky130_fd_sc_hd__dfrtp_2 _5245_ (.CLK(clk),
    .D(_0425_),
    .RESET_B(_1144_),
    .Q(\gen_pe[3].pe_inst.out_right[17] ));
 sky130_fd_sc_hd__dfrtp_2 _5246_ (.CLK(clk),
    .D(_0426_),
    .RESET_B(_1145_),
    .Q(\gen_pe[3].pe_inst.out_right[18] ));
 sky130_fd_sc_hd__dfrtp_2 _5247_ (.CLK(clk),
    .D(_0427_),
    .RESET_B(_1146_),
    .Q(\gen_pe[3].pe_inst.out_right[19] ));
 sky130_fd_sc_hd__dfrtp_2 _5248_ (.CLK(clk),
    .D(_0429_),
    .RESET_B(_1147_),
    .Q(\gen_pe[3].pe_inst.out_right[20] ));
 sky130_fd_sc_hd__dfrtp_2 _5249_ (.CLK(clk),
    .D(_0430_),
    .RESET_B(_1148_),
    .Q(\gen_pe[3].pe_inst.out_right[21] ));
 sky130_fd_sc_hd__dfrtp_2 _5250_ (.CLK(clk),
    .D(_0431_),
    .RESET_B(_1149_),
    .Q(\gen_pe[3].pe_inst.out_right[22] ));
 sky130_fd_sc_hd__dfrtp_2 _5251_ (.CLK(clk),
    .D(_0432_),
    .RESET_B(_1150_),
    .Q(\gen_pe[3].pe_inst.out_right[23] ));
 sky130_fd_sc_hd__dfrtp_2 _5252_ (.CLK(clk),
    .D(_0433_),
    .RESET_B(_1151_),
    .Q(\gen_pe[3].pe_inst.out_right[24] ));
 sky130_fd_sc_hd__dfrtp_2 _5253_ (.CLK(clk),
    .D(_0434_),
    .RESET_B(_1152_),
    .Q(\gen_pe[3].pe_inst.out_right[25] ));
 sky130_fd_sc_hd__dfrtp_2 _5254_ (.CLK(clk),
    .D(_0435_),
    .RESET_B(_1153_),
    .Q(\gen_pe[3].pe_inst.out_right[26] ));
 sky130_fd_sc_hd__dfrtp_2 _5255_ (.CLK(clk),
    .D(_0436_),
    .RESET_B(_1154_),
    .Q(\gen_pe[3].pe_inst.out_right[27] ));
 sky130_fd_sc_hd__dfrtp_2 _5256_ (.CLK(clk),
    .D(_0437_),
    .RESET_B(_1155_),
    .Q(\gen_pe[3].pe_inst.out_right[28] ));
 sky130_fd_sc_hd__dfrtp_2 _5257_ (.CLK(clk),
    .D(_0438_),
    .RESET_B(_1156_),
    .Q(\gen_pe[3].pe_inst.out_right[29] ));
 sky130_fd_sc_hd__dfrtp_2 _5258_ (.CLK(clk),
    .D(_0440_),
    .RESET_B(_1157_),
    .Q(\gen_pe[3].pe_inst.out_right[30] ));
 sky130_fd_sc_hd__dfrtp_2 _5259_ (.CLK(clk),
    .D(_0441_),
    .RESET_B(_1158_),
    .Q(\gen_pe[3].pe_inst.out_right[31] ));
 sky130_fd_sc_hd__dfrtp_2 _5260_ (.CLK(clk),
    .D(_0577_),
    .RESET_B(_1159_),
    .Q(\gen_left[6][0] ));
 sky130_fd_sc_hd__dfrtp_2 _5261_ (.CLK(clk),
    .D(_0588_),
    .RESET_B(_1160_),
    .Q(\gen_left[6][1] ));
 sky130_fd_sc_hd__dfrtp_2 _5262_ (.CLK(clk),
    .D(_0599_),
    .RESET_B(_1161_),
    .Q(\gen_left[6][2] ));
 sky130_fd_sc_hd__dfrtp_2 _5263_ (.CLK(clk),
    .D(_0602_),
    .RESET_B(_1162_),
    .Q(\gen_left[6][3] ));
 sky130_fd_sc_hd__dfrtp_2 _5264_ (.CLK(clk),
    .D(_0603_),
    .RESET_B(_1163_),
    .Q(\gen_left[6][4] ));
 sky130_fd_sc_hd__dfrtp_2 _5265_ (.CLK(clk),
    .D(_0604_),
    .RESET_B(_1164_),
    .Q(\gen_left[6][5] ));
 sky130_fd_sc_hd__dfrtp_2 _5266_ (.CLK(clk),
    .D(_0605_),
    .RESET_B(_1165_),
    .Q(\gen_left[6][6] ));
 sky130_fd_sc_hd__dfrtp_2 _5267_ (.CLK(clk),
    .D(_0606_),
    .RESET_B(_1166_),
    .Q(\gen_left[6][7] ));
 sky130_fd_sc_hd__dfrtp_2 _5268_ (.CLK(clk),
    .D(_0607_),
    .RESET_B(_1167_),
    .Q(\gen_left[6][8] ));
 sky130_fd_sc_hd__dfrtp_2 _5269_ (.CLK(clk),
    .D(_0608_),
    .RESET_B(_1168_),
    .Q(\gen_left[6][9] ));
 sky130_fd_sc_hd__dfrtp_2 _5270_ (.CLK(clk),
    .D(_0578_),
    .RESET_B(_1169_),
    .Q(\gen_left[6][10] ));
 sky130_fd_sc_hd__dfrtp_2 _5271_ (.CLK(clk),
    .D(_0579_),
    .RESET_B(_1170_),
    .Q(\gen_left[6][11] ));
 sky130_fd_sc_hd__dfrtp_2 _5272_ (.CLK(clk),
    .D(_0580_),
    .RESET_B(_1171_),
    .Q(\gen_left[6][12] ));
 sky130_fd_sc_hd__dfrtp_2 _5273_ (.CLK(clk),
    .D(_0581_),
    .RESET_B(_1172_),
    .Q(\gen_left[6][13] ));
 sky130_fd_sc_hd__dfrtp_2 _5274_ (.CLK(clk),
    .D(_0582_),
    .RESET_B(_1173_),
    .Q(\gen_left[6][14] ));
 sky130_fd_sc_hd__dfrtp_2 _5275_ (.CLK(clk),
    .D(_0583_),
    .RESET_B(_1174_),
    .Q(\gen_left[6][15] ));
 sky130_fd_sc_hd__dfrtp_2 _5276_ (.CLK(clk),
    .D(_0584_),
    .RESET_B(_1175_),
    .Q(\gen_left[6][16] ));
 sky130_fd_sc_hd__dfrtp_2 _5277_ (.CLK(clk),
    .D(_0585_),
    .RESET_B(_1176_),
    .Q(\gen_left[6][17] ));
 sky130_fd_sc_hd__dfrtp_2 _5278_ (.CLK(clk),
    .D(_0586_),
    .RESET_B(_1177_),
    .Q(\gen_left[6][18] ));
 sky130_fd_sc_hd__dfrtp_2 _5279_ (.CLK(clk),
    .D(_0587_),
    .RESET_B(_1178_),
    .Q(\gen_left[6][19] ));
 sky130_fd_sc_hd__dfrtp_2 _5280_ (.CLK(clk),
    .D(_0589_),
    .RESET_B(_1179_),
    .Q(\gen_left[6][20] ));
 sky130_fd_sc_hd__dfrtp_2 _5281_ (.CLK(clk),
    .D(_0590_),
    .RESET_B(_1180_),
    .Q(\gen_left[6][21] ));
 sky130_fd_sc_hd__dfrtp_2 _5282_ (.CLK(clk),
    .D(_0591_),
    .RESET_B(_1181_),
    .Q(\gen_left[6][22] ));
 sky130_fd_sc_hd__dfrtp_2 _5283_ (.CLK(clk),
    .D(_0592_),
    .RESET_B(_1182_),
    .Q(\gen_left[6][23] ));
 sky130_fd_sc_hd__dfrtp_2 _5284_ (.CLK(clk),
    .D(_0593_),
    .RESET_B(_1183_),
    .Q(\gen_left[6][24] ));
 sky130_fd_sc_hd__dfrtp_2 _5285_ (.CLK(clk),
    .D(_0594_),
    .RESET_B(_1184_),
    .Q(\gen_left[6][25] ));
 sky130_fd_sc_hd__dfrtp_2 _5286_ (.CLK(clk),
    .D(_0595_),
    .RESET_B(_1185_),
    .Q(\gen_left[6][26] ));
 sky130_fd_sc_hd__dfrtp_2 _5287_ (.CLK(clk),
    .D(_0596_),
    .RESET_B(_1186_),
    .Q(\gen_left[6][27] ));
 sky130_fd_sc_hd__dfrtp_2 _5288_ (.CLK(clk),
    .D(_0597_),
    .RESET_B(_1187_),
    .Q(\gen_left[6][28] ));
 sky130_fd_sc_hd__dfrtp_2 _5289_ (.CLK(clk),
    .D(_0598_),
    .RESET_B(_1188_),
    .Q(\gen_left[6][29] ));
 sky130_fd_sc_hd__dfrtp_2 _5290_ (.CLK(clk),
    .D(_0600_),
    .RESET_B(_1189_),
    .Q(\gen_left[6][30] ));
 sky130_fd_sc_hd__dfrtp_2 _5291_ (.CLK(clk),
    .D(_0601_),
    .RESET_B(_1190_),
    .Q(\gen_left[6][31] ));
 sky130_fd_sc_hd__dfrtp_2 _5292_ (.CLK(clk),
    .D(_1346_),
    .RESET_B(_1191_),
    .Q(out_data_flat[224]));
 sky130_fd_sc_hd__dfrtp_2 _5293_ (.CLK(clk),
    .D(_1347_),
    .RESET_B(_1192_),
    .Q(out_data_flat[225]));
 sky130_fd_sc_hd__dfrtp_2 _5294_ (.CLK(clk),
    .D(_1348_),
    .RESET_B(_1193_),
    .Q(out_data_flat[226]));
 sky130_fd_sc_hd__dfrtp_2 _5295_ (.CLK(clk),
    .D(_1349_),
    .RESET_B(_1194_),
    .Q(out_data_flat[227]));
 sky130_fd_sc_hd__dfrtp_2 _5296_ (.CLK(clk),
    .D(_1350_),
    .RESET_B(_1195_),
    .Q(out_data_flat[228]));
 sky130_fd_sc_hd__dfrtp_2 _5297_ (.CLK(clk),
    .D(_1351_),
    .RESET_B(_1196_),
    .Q(out_data_flat[229]));
 sky130_fd_sc_hd__dfrtp_2 _5298_ (.CLK(clk),
    .D(_1352_),
    .RESET_B(_1197_),
    .Q(out_data_flat[230]));
 sky130_fd_sc_hd__dfrtp_2 _5299_ (.CLK(clk),
    .D(_1353_),
    .RESET_B(_1198_),
    .Q(out_data_flat[231]));
 sky130_fd_sc_hd__dfrtp_2 _5300_ (.CLK(clk),
    .D(_1354_),
    .RESET_B(_1199_),
    .Q(out_data_flat[232]));
 sky130_fd_sc_hd__dfrtp_2 _5301_ (.CLK(clk),
    .D(_1355_),
    .RESET_B(_1200_),
    .Q(out_data_flat[233]));
 sky130_fd_sc_hd__dfrtp_2 _5302_ (.CLK(clk),
    .D(_1356_),
    .RESET_B(_1201_),
    .Q(out_data_flat[234]));
 sky130_fd_sc_hd__dfrtp_2 _5303_ (.CLK(clk),
    .D(_1357_),
    .RESET_B(_1202_),
    .Q(out_data_flat[235]));
 sky130_fd_sc_hd__dfrtp_2 _5304_ (.CLK(clk),
    .D(_1358_),
    .RESET_B(_1203_),
    .Q(out_data_flat[236]));
 sky130_fd_sc_hd__dfrtp_2 _5305_ (.CLK(clk),
    .D(_1359_),
    .RESET_B(_1204_),
    .Q(out_data_flat[237]));
 sky130_fd_sc_hd__dfrtp_2 _5306_ (.CLK(clk),
    .D(_1360_),
    .RESET_B(_1205_),
    .Q(out_data_flat[238]));
 sky130_fd_sc_hd__dfrtp_2 _5307_ (.CLK(clk),
    .D(_1361_),
    .RESET_B(_1206_),
    .Q(out_data_flat[239]));
 sky130_fd_sc_hd__dfrtp_2 _5308_ (.CLK(clk),
    .D(_1362_),
    .RESET_B(_1207_),
    .Q(out_data_flat[240]));
 sky130_fd_sc_hd__dfrtp_2 _5309_ (.CLK(clk),
    .D(_1363_),
    .RESET_B(_1208_),
    .Q(out_data_flat[241]));
 sky130_fd_sc_hd__dfrtp_2 _5310_ (.CLK(clk),
    .D(_1364_),
    .RESET_B(_1209_),
    .Q(out_data_flat[242]));
 sky130_fd_sc_hd__dfrtp_2 _5311_ (.CLK(clk),
    .D(_1365_),
    .RESET_B(_1210_),
    .Q(out_data_flat[243]));
 sky130_fd_sc_hd__dfrtp_2 _5312_ (.CLK(clk),
    .D(_1366_),
    .RESET_B(_1211_),
    .Q(out_data_flat[244]));
 sky130_fd_sc_hd__dfrtp_2 _5313_ (.CLK(clk),
    .D(_1367_),
    .RESET_B(_1212_),
    .Q(out_data_flat[245]));
 sky130_fd_sc_hd__dfrtp_2 _5314_ (.CLK(clk),
    .D(_1368_),
    .RESET_B(_1213_),
    .Q(out_data_flat[246]));
 sky130_fd_sc_hd__dfrtp_2 _5315_ (.CLK(clk),
    .D(_1369_),
    .RESET_B(_1214_),
    .Q(out_data_flat[247]));
 sky130_fd_sc_hd__dfrtp_2 _5316_ (.CLK(clk),
    .D(_1370_),
    .RESET_B(_1215_),
    .Q(out_data_flat[248]));
 sky130_fd_sc_hd__dfrtp_2 _5317_ (.CLK(clk),
    .D(_1371_),
    .RESET_B(_1216_),
    .Q(out_data_flat[249]));
 sky130_fd_sc_hd__dfrtp_2 _5318_ (.CLK(clk),
    .D(_1372_),
    .RESET_B(_1217_),
    .Q(out_data_flat[250]));
 sky130_fd_sc_hd__dfrtp_2 _5319_ (.CLK(clk),
    .D(_1373_),
    .RESET_B(_1218_),
    .Q(out_data_flat[251]));
 sky130_fd_sc_hd__dfrtp_2 _5320_ (.CLK(clk),
    .D(_1374_),
    .RESET_B(_1219_),
    .Q(out_data_flat[252]));
 sky130_fd_sc_hd__dfrtp_2 _5321_ (.CLK(clk),
    .D(_1375_),
    .RESET_B(_1220_),
    .Q(out_data_flat[253]));
 sky130_fd_sc_hd__dfrtp_2 _5322_ (.CLK(clk),
    .D(_1376_),
    .RESET_B(_1221_),
    .Q(out_data_flat[254]));
 sky130_fd_sc_hd__dfrtp_2 _5323_ (.CLK(clk),
    .D(_1377_),
    .RESET_B(_1222_),
    .Q(out_data_flat[255]));
 sky130_fd_sc_hd__dfrtp_2 _5324_ (.CLK(clk),
    .D(_1378_),
    .RESET_B(_1223_),
    .Q(out_data_flat[0]));
 sky130_fd_sc_hd__dfrtp_2 _5325_ (.CLK(clk),
    .D(_1379_),
    .RESET_B(_1224_),
    .Q(out_data_flat[1]));
 sky130_fd_sc_hd__dfrtp_2 _5326_ (.CLK(clk),
    .D(_1380_),
    .RESET_B(_1225_),
    .Q(out_data_flat[2]));
 sky130_fd_sc_hd__dfrtp_2 _5327_ (.CLK(clk),
    .D(_1381_),
    .RESET_B(_1226_),
    .Q(out_data_flat[3]));
 sky130_fd_sc_hd__dfrtp_2 _5328_ (.CLK(clk),
    .D(_1382_),
    .RESET_B(_1227_),
    .Q(out_data_flat[4]));
 sky130_fd_sc_hd__dfrtp_2 _5329_ (.CLK(clk),
    .D(_1383_),
    .RESET_B(_1228_),
    .Q(out_data_flat[5]));
 sky130_fd_sc_hd__dfrtp_2 _5330_ (.CLK(clk),
    .D(_1384_),
    .RESET_B(_1229_),
    .Q(out_data_flat[6]));
 sky130_fd_sc_hd__dfrtp_2 _5331_ (.CLK(clk),
    .D(_1385_),
    .RESET_B(_1230_),
    .Q(out_data_flat[7]));
 sky130_fd_sc_hd__dfrtp_2 _5332_ (.CLK(clk),
    .D(_1386_),
    .RESET_B(_1231_),
    .Q(out_data_flat[8]));
 sky130_fd_sc_hd__dfrtp_2 _5333_ (.CLK(clk),
    .D(_1387_),
    .RESET_B(_1232_),
    .Q(out_data_flat[9]));
 sky130_fd_sc_hd__dfrtp_2 _5334_ (.CLK(clk),
    .D(_1388_),
    .RESET_B(_1233_),
    .Q(out_data_flat[10]));
 sky130_fd_sc_hd__dfrtp_2 _5335_ (.CLK(clk),
    .D(_1389_),
    .RESET_B(_1234_),
    .Q(out_data_flat[11]));
 sky130_fd_sc_hd__dfrtp_2 _5336_ (.CLK(clk),
    .D(_1390_),
    .RESET_B(_1235_),
    .Q(out_data_flat[12]));
 sky130_fd_sc_hd__dfrtp_2 _5337_ (.CLK(clk),
    .D(_1391_),
    .RESET_B(_1236_),
    .Q(out_data_flat[13]));
 sky130_fd_sc_hd__dfrtp_2 _5338_ (.CLK(clk),
    .D(_1392_),
    .RESET_B(_1237_),
    .Q(out_data_flat[14]));
 sky130_fd_sc_hd__dfrtp_2 _5339_ (.CLK(clk),
    .D(_1393_),
    .RESET_B(_1238_),
    .Q(out_data_flat[15]));
 sky130_fd_sc_hd__dfrtp_2 _5340_ (.CLK(clk),
    .D(_1394_),
    .RESET_B(_1239_),
    .Q(out_data_flat[16]));
 sky130_fd_sc_hd__dfrtp_2 _5341_ (.CLK(clk),
    .D(_1395_),
    .RESET_B(_1240_),
    .Q(out_data_flat[17]));
 sky130_fd_sc_hd__dfrtp_2 _5342_ (.CLK(clk),
    .D(_1396_),
    .RESET_B(_1241_),
    .Q(out_data_flat[18]));
 sky130_fd_sc_hd__dfrtp_2 _5343_ (.CLK(clk),
    .D(_1397_),
    .RESET_B(_1242_),
    .Q(out_data_flat[19]));
 sky130_fd_sc_hd__dfrtp_2 _5344_ (.CLK(clk),
    .D(_1398_),
    .RESET_B(_1243_),
    .Q(out_data_flat[20]));
 sky130_fd_sc_hd__dfrtp_2 _5345_ (.CLK(clk),
    .D(_1399_),
    .RESET_B(_1244_),
    .Q(out_data_flat[21]));
 sky130_fd_sc_hd__dfrtp_2 _5346_ (.CLK(clk),
    .D(_1400_),
    .RESET_B(_1245_),
    .Q(out_data_flat[22]));
 sky130_fd_sc_hd__dfrtp_2 _5347_ (.CLK(clk),
    .D(_1401_),
    .RESET_B(_1246_),
    .Q(out_data_flat[23]));
 sky130_fd_sc_hd__dfrtp_2 _5348_ (.CLK(clk),
    .D(_1402_),
    .RESET_B(_1247_),
    .Q(out_data_flat[24]));
 sky130_fd_sc_hd__dfrtp_2 _5349_ (.CLK(clk),
    .D(_1403_),
    .RESET_B(_1248_),
    .Q(out_data_flat[25]));
 sky130_fd_sc_hd__dfrtp_2 _5350_ (.CLK(clk),
    .D(_1404_),
    .RESET_B(_1249_),
    .Q(out_data_flat[26]));
 sky130_fd_sc_hd__dfrtp_2 _5351_ (.CLK(clk),
    .D(_1405_),
    .RESET_B(_1250_),
    .Q(out_data_flat[27]));
 sky130_fd_sc_hd__dfrtp_2 _5352_ (.CLK(clk),
    .D(_1406_),
    .RESET_B(_1251_),
    .Q(out_data_flat[28]));
 sky130_fd_sc_hd__dfrtp_2 _5353_ (.CLK(clk),
    .D(_1407_),
    .RESET_B(_1252_),
    .Q(out_data_flat[29]));
 sky130_fd_sc_hd__dfrtp_2 _5354_ (.CLK(clk),
    .D(_1408_),
    .RESET_B(_1253_),
    .Q(out_data_flat[30]));
 sky130_fd_sc_hd__dfrtp_2 _5355_ (.CLK(clk),
    .D(_1409_),
    .RESET_B(_1254_),
    .Q(out_data_flat[31]));
 sky130_fd_sc_hd__dfrtp_2 _5356_ (.CLK(clk),
    .D(_0160_),
    .RESET_B(_1255_),
    .Q(out_data_flat[192]));
 sky130_fd_sc_hd__dfrtp_2 _5357_ (.CLK(clk),
    .D(_0171_),
    .RESET_B(_1256_),
    .Q(out_data_flat[193]));
 sky130_fd_sc_hd__dfrtp_2 _5358_ (.CLK(clk),
    .D(_0182_),
    .RESET_B(_1257_),
    .Q(out_data_flat[194]));
 sky130_fd_sc_hd__dfrtp_2 _5359_ (.CLK(clk),
    .D(_0185_),
    .RESET_B(_1258_),
    .Q(out_data_flat[195]));
 sky130_fd_sc_hd__dfrtp_2 _5360_ (.CLK(clk),
    .D(_0186_),
    .RESET_B(_1259_),
    .Q(out_data_flat[196]));
 sky130_fd_sc_hd__dfrtp_2 _5361_ (.CLK(clk),
    .D(_0187_),
    .RESET_B(_1260_),
    .Q(out_data_flat[197]));
 sky130_fd_sc_hd__dfrtp_2 _5362_ (.CLK(clk),
    .D(_0188_),
    .RESET_B(_1261_),
    .Q(out_data_flat[198]));
 sky130_fd_sc_hd__dfrtp_2 _5363_ (.CLK(clk),
    .D(_0189_),
    .RESET_B(_1262_),
    .Q(out_data_flat[199]));
 sky130_fd_sc_hd__dfrtp_2 _5364_ (.CLK(clk),
    .D(_0190_),
    .RESET_B(_1263_),
    .Q(out_data_flat[200]));
 sky130_fd_sc_hd__dfrtp_2 _5365_ (.CLK(clk),
    .D(_0191_),
    .RESET_B(_1264_),
    .Q(out_data_flat[201]));
 sky130_fd_sc_hd__dfrtp_2 _5366_ (.CLK(clk),
    .D(_0161_),
    .RESET_B(_1265_),
    .Q(out_data_flat[202]));
 sky130_fd_sc_hd__dfrtp_2 _5367_ (.CLK(clk),
    .D(_0162_),
    .RESET_B(_1266_),
    .Q(out_data_flat[203]));
 sky130_fd_sc_hd__dfrtp_2 _5368_ (.CLK(clk),
    .D(_0163_),
    .RESET_B(_1267_),
    .Q(out_data_flat[204]));
 sky130_fd_sc_hd__dfrtp_2 _5369_ (.CLK(clk),
    .D(_0164_),
    .RESET_B(_1268_),
    .Q(out_data_flat[205]));
 sky130_fd_sc_hd__dfrtp_2 _5370_ (.CLK(clk),
    .D(_0165_),
    .RESET_B(_1269_),
    .Q(out_data_flat[206]));
 sky130_fd_sc_hd__dfrtp_2 _5371_ (.CLK(clk),
    .D(_0166_),
    .RESET_B(_1270_),
    .Q(out_data_flat[207]));
 sky130_fd_sc_hd__dfrtp_2 _5372_ (.CLK(clk),
    .D(_0167_),
    .RESET_B(_1271_),
    .Q(out_data_flat[208]));
 sky130_fd_sc_hd__dfrtp_2 _5373_ (.CLK(clk),
    .D(_0168_),
    .RESET_B(_1272_),
    .Q(out_data_flat[209]));
 sky130_fd_sc_hd__dfrtp_2 _5374_ (.CLK(clk),
    .D(_0169_),
    .RESET_B(_1273_),
    .Q(out_data_flat[210]));
 sky130_fd_sc_hd__dfrtp_2 _5375_ (.CLK(clk),
    .D(_0170_),
    .RESET_B(_1274_),
    .Q(out_data_flat[211]));
 sky130_fd_sc_hd__dfrtp_2 _5376_ (.CLK(clk),
    .D(_0172_),
    .RESET_B(_1275_),
    .Q(out_data_flat[212]));
 sky130_fd_sc_hd__dfrtp_2 _5377_ (.CLK(clk),
    .D(_0173_),
    .RESET_B(_1276_),
    .Q(out_data_flat[213]));
 sky130_fd_sc_hd__dfrtp_2 _5378_ (.CLK(clk),
    .D(_0174_),
    .RESET_B(_1277_),
    .Q(out_data_flat[214]));
 sky130_fd_sc_hd__dfrtp_2 _5379_ (.CLK(clk),
    .D(_0175_),
    .RESET_B(_1278_),
    .Q(out_data_flat[215]));
 sky130_fd_sc_hd__dfrtp_2 _5380_ (.CLK(clk),
    .D(_0176_),
    .RESET_B(_1279_),
    .Q(out_data_flat[216]));
 sky130_fd_sc_hd__dfrtp_2 _5381_ (.CLK(clk),
    .D(_0177_),
    .RESET_B(_1280_),
    .Q(out_data_flat[217]));
 sky130_fd_sc_hd__dfrtp_2 _5382_ (.CLK(clk),
    .D(_0178_),
    .RESET_B(_1281_),
    .Q(out_data_flat[218]));
 sky130_fd_sc_hd__dfrtp_2 _5383_ (.CLK(clk),
    .D(_0179_),
    .RESET_B(_1282_),
    .Q(out_data_flat[219]));
 sky130_fd_sc_hd__dfrtp_2 _5384_ (.CLK(clk),
    .D(_0180_),
    .RESET_B(_1283_),
    .Q(out_data_flat[220]));
 sky130_fd_sc_hd__dfrtp_2 _5385_ (.CLK(clk),
    .D(_0181_),
    .RESET_B(_1284_),
    .Q(out_data_flat[221]));
 sky130_fd_sc_hd__dfrtp_2 _5386_ (.CLK(clk),
    .D(_0183_),
    .RESET_B(_1285_),
    .Q(out_data_flat[222]));
 sky130_fd_sc_hd__dfrtp_2 _5387_ (.CLK(clk),
    .D(_0184_),
    .RESET_B(_1286_),
    .Q(out_data_flat[223]));
 sky130_fd_sc_hd__dfrtp_2 _5388_ (.CLK(clk),
    .D(_0128_),
    .RESET_B(_1287_),
    .Q(out_data_flat[160]));
 sky130_fd_sc_hd__dfrtp_2 _5389_ (.CLK(clk),
    .D(_0139_),
    .RESET_B(_1288_),
    .Q(out_data_flat[161]));
 sky130_fd_sc_hd__dfrtp_2 _5390_ (.CLK(clk),
    .D(_0150_),
    .RESET_B(_1289_),
    .Q(out_data_flat[162]));
 sky130_fd_sc_hd__dfrtp_2 _5391_ (.CLK(clk),
    .D(_0153_),
    .RESET_B(_1290_),
    .Q(out_data_flat[163]));
 sky130_fd_sc_hd__dfrtp_2 _5392_ (.CLK(clk),
    .D(_0154_),
    .RESET_B(_1291_),
    .Q(out_data_flat[164]));
 sky130_fd_sc_hd__dfrtp_2 _5393_ (.CLK(clk),
    .D(_0155_),
    .RESET_B(_1292_),
    .Q(out_data_flat[165]));
 sky130_fd_sc_hd__dfrtp_2 _5394_ (.CLK(clk),
    .D(_0156_),
    .RESET_B(_1293_),
    .Q(out_data_flat[166]));
 sky130_fd_sc_hd__dfrtp_2 _5395_ (.CLK(clk),
    .D(_0157_),
    .RESET_B(_1294_),
    .Q(out_data_flat[167]));
 sky130_fd_sc_hd__dfrtp_2 _5396_ (.CLK(clk),
    .D(_0158_),
    .RESET_B(_1295_),
    .Q(out_data_flat[168]));
 sky130_fd_sc_hd__dfrtp_2 _5397_ (.CLK(clk),
    .D(_0159_),
    .RESET_B(_1296_),
    .Q(out_data_flat[169]));
 sky130_fd_sc_hd__dfrtp_2 _5398_ (.CLK(clk),
    .D(_0129_),
    .RESET_B(_1297_),
    .Q(out_data_flat[170]));
 sky130_fd_sc_hd__dfrtp_2 _5399_ (.CLK(clk),
    .D(_0130_),
    .RESET_B(_1298_),
    .Q(out_data_flat[171]));
 sky130_fd_sc_hd__dfrtp_2 _5400_ (.CLK(clk),
    .D(_0131_),
    .RESET_B(_1299_),
    .Q(out_data_flat[172]));
 sky130_fd_sc_hd__dfrtp_2 _5401_ (.CLK(clk),
    .D(_0132_),
    .RESET_B(_1300_),
    .Q(out_data_flat[173]));
 sky130_fd_sc_hd__dfrtp_2 _5402_ (.CLK(clk),
    .D(_0133_),
    .RESET_B(_1301_),
    .Q(out_data_flat[174]));
 sky130_fd_sc_hd__dfrtp_2 _5403_ (.CLK(clk),
    .D(_0134_),
    .RESET_B(_1302_),
    .Q(out_data_flat[175]));
 sky130_fd_sc_hd__dfrtp_2 _5404_ (.CLK(clk),
    .D(_0135_),
    .RESET_B(_1303_),
    .Q(out_data_flat[176]));
 sky130_fd_sc_hd__dfrtp_2 _5405_ (.CLK(clk),
    .D(_0136_),
    .RESET_B(_1304_),
    .Q(out_data_flat[177]));
 sky130_fd_sc_hd__dfrtp_2 _5406_ (.CLK(clk),
    .D(_0137_),
    .RESET_B(_1305_),
    .Q(out_data_flat[178]));
 sky130_fd_sc_hd__dfrtp_2 _5407_ (.CLK(clk),
    .D(_0138_),
    .RESET_B(_1306_),
    .Q(out_data_flat[179]));
 sky130_fd_sc_hd__dfrtp_2 _5408_ (.CLK(clk),
    .D(_0140_),
    .RESET_B(_1307_),
    .Q(out_data_flat[180]));
 sky130_fd_sc_hd__dfrtp_2 _5409_ (.CLK(clk),
    .D(_0141_),
    .RESET_B(_1308_),
    .Q(out_data_flat[181]));
 sky130_fd_sc_hd__dfrtp_2 _5410_ (.CLK(clk),
    .D(_0142_),
    .RESET_B(_1309_),
    .Q(out_data_flat[182]));
 sky130_fd_sc_hd__dfrtp_2 _5411_ (.CLK(clk),
    .D(_0143_),
    .RESET_B(_1310_),
    .Q(out_data_flat[183]));
 sky130_fd_sc_hd__dfrtp_2 _5412_ (.CLK(clk),
    .D(_0144_),
    .RESET_B(_1311_),
    .Q(out_data_flat[184]));
 sky130_fd_sc_hd__dfrtp_2 _5413_ (.CLK(clk),
    .D(_0145_),
    .RESET_B(_1312_),
    .Q(out_data_flat[185]));
 sky130_fd_sc_hd__dfrtp_2 _5414_ (.CLK(clk),
    .D(_0146_),
    .RESET_B(_1313_),
    .Q(out_data_flat[186]));
 sky130_fd_sc_hd__dfrtp_2 _5415_ (.CLK(clk),
    .D(_0147_),
    .RESET_B(_1314_),
    .Q(out_data_flat[187]));
 sky130_fd_sc_hd__dfrtp_2 _5416_ (.CLK(clk),
    .D(_0148_),
    .RESET_B(_1315_),
    .Q(out_data_flat[188]));
 sky130_fd_sc_hd__dfrtp_2 _5417_ (.CLK(clk),
    .D(_0149_),
    .RESET_B(_1316_),
    .Q(out_data_flat[189]));
 sky130_fd_sc_hd__dfrtp_2 _5418_ (.CLK(clk),
    .D(_0151_),
    .RESET_B(_1317_),
    .Q(out_data_flat[190]));
 sky130_fd_sc_hd__dfrtp_2 _5419_ (.CLK(clk),
    .D(_0152_),
    .RESET_B(_1318_),
    .Q(out_data_flat[191]));
 sky130_fd_sc_hd__dfrtp_2 _5420_ (.CLK(clk),
    .D(_0096_),
    .RESET_B(_1319_),
    .Q(out_data_flat[128]));
 sky130_fd_sc_hd__dfrtp_2 _5421_ (.CLK(clk),
    .D(_0107_),
    .RESET_B(_1320_),
    .Q(out_data_flat[129]));
 sky130_fd_sc_hd__dfrtp_2 _5422_ (.CLK(clk),
    .D(_0118_),
    .RESET_B(_1321_),
    .Q(out_data_flat[130]));
 sky130_fd_sc_hd__dfrtp_2 _5423_ (.CLK(clk),
    .D(_0121_),
    .RESET_B(_1322_),
    .Q(out_data_flat[131]));
 sky130_fd_sc_hd__dfrtp_2 _5424_ (.CLK(clk),
    .D(_0122_),
    .RESET_B(_1323_),
    .Q(out_data_flat[132]));
 sky130_fd_sc_hd__dfrtp_2 _5425_ (.CLK(clk),
    .D(_0123_),
    .RESET_B(_1324_),
    .Q(out_data_flat[133]));
 sky130_fd_sc_hd__dfrtp_2 _5426_ (.CLK(clk),
    .D(_0124_),
    .RESET_B(_1325_),
    .Q(out_data_flat[134]));
 sky130_fd_sc_hd__dfrtp_2 _5427_ (.CLK(clk),
    .D(_0125_),
    .RESET_B(_1326_),
    .Q(out_data_flat[135]));
 sky130_fd_sc_hd__dfrtp_2 _5428_ (.CLK(clk),
    .D(_0126_),
    .RESET_B(_1327_),
    .Q(out_data_flat[136]));
 sky130_fd_sc_hd__dfrtp_2 _5429_ (.CLK(clk),
    .D(_0127_),
    .RESET_B(_1328_),
    .Q(out_data_flat[137]));
 sky130_fd_sc_hd__dfrtp_2 _5430_ (.CLK(clk),
    .D(_0097_),
    .RESET_B(_1329_),
    .Q(out_data_flat[138]));
 sky130_fd_sc_hd__dfrtp_2 _5431_ (.CLK(clk),
    .D(_0098_),
    .RESET_B(_1330_),
    .Q(out_data_flat[139]));
 sky130_fd_sc_hd__dfrtp_2 _5432_ (.CLK(clk),
    .D(_0099_),
    .RESET_B(_1331_),
    .Q(out_data_flat[140]));
 sky130_fd_sc_hd__dfrtp_2 _5433_ (.CLK(clk),
    .D(_0100_),
    .RESET_B(_1332_),
    .Q(out_data_flat[141]));
 sky130_fd_sc_hd__dfrtp_2 _5434_ (.CLK(clk),
    .D(_0101_),
    .RESET_B(_1333_),
    .Q(out_data_flat[142]));
 sky130_fd_sc_hd__dfrtp_2 _5435_ (.CLK(clk),
    .D(_0102_),
    .RESET_B(_1334_),
    .Q(out_data_flat[143]));
 sky130_fd_sc_hd__dfrtp_2 _5436_ (.CLK(clk),
    .D(_0103_),
    .RESET_B(_1335_),
    .Q(out_data_flat[144]));
 sky130_fd_sc_hd__dfrtp_2 _5437_ (.CLK(clk),
    .D(_0104_),
    .RESET_B(_1336_),
    .Q(out_data_flat[145]));
 sky130_fd_sc_hd__dfrtp_2 _5438_ (.CLK(clk),
    .D(_0105_),
    .RESET_B(_1337_),
    .Q(out_data_flat[146]));
 sky130_fd_sc_hd__dfrtp_2 _5439_ (.CLK(clk),
    .D(_0106_),
    .RESET_B(_1338_),
    .Q(out_data_flat[147]));
 sky130_fd_sc_hd__dfrtp_2 _5440_ (.CLK(clk),
    .D(_0108_),
    .RESET_B(_1339_),
    .Q(out_data_flat[148]));
 sky130_fd_sc_hd__dfrtp_2 _5441_ (.CLK(clk),
    .D(_0109_),
    .RESET_B(_1340_),
    .Q(out_data_flat[149]));
 sky130_fd_sc_hd__dfrtp_2 _5442_ (.CLK(clk),
    .D(_0110_),
    .RESET_B(_1341_),
    .Q(out_data_flat[150]));
 sky130_fd_sc_hd__dfrtp_2 _5443_ (.CLK(clk),
    .D(_0111_),
    .RESET_B(_1342_),
    .Q(out_data_flat[151]));
 sky130_fd_sc_hd__dfrtp_2 _5444_ (.CLK(clk),
    .D(_0112_),
    .RESET_B(_1343_),
    .Q(out_data_flat[152]));
 sky130_fd_sc_hd__dfrtp_2 _5445_ (.CLK(clk),
    .D(_0113_),
    .RESET_B(_1344_),
    .Q(out_data_flat[153]));
 sky130_fd_sc_hd__dfrtp_2 _5446_ (.CLK(clk),
    .D(_0114_),
    .RESET_B(_1345_),
    .Q(out_data_flat[154]));
endmodule
