`timescale 1ns / 1ps

module mac4_tb;

    logic signed [15:0] a0, b0;
    logic signed [15:0] a1, b1;
    logic signed [15:0] a2, b2;
    logic signed [15:0] a3, b3;
    logic signed [15:0] result;

    // Instantiate DUT
    mac4 dut (
        .a0(a0), .b0(b0),
        .a1(a1), .b1(b1),
        .a2(a2), .b2(b2),
        .a3(a3), .b3(b3),
        .result(result)
    );

    initial begin
        // Test case 1
        // Each product will be: (Q2.14 * Q4.12) = Q6.26 → >>>14 → Q4.12
        //
        // a0 = 0.5  (Q2.14) =  0b_0010_0000_0000_0000 = 8192
        // b0 = 2.0  (Q4.12) =  0b_0010_0000_0000_0000 = 8192
        // a1 = 1.0  (Q2.14) =  0b_0100_0000_0000_0000 = 16384
        // b1 = 1.0  (Q4.12) =  0b_0001_0000_0000_0000 = 4096
        // a2 = -0.5 (Q2.14) =  0b_1110_0000_0000_0000 = -8192
        // b2 = 1.0  (Q4.12) =  0b_0001_0000_0000_0000 = 4096
        // a3 = 0.25 (Q2.14) =  0b_0001_0000_0000_0000 = 4096
        // b3 = 4.0  (Q4.12) =  0b_0100_0000_0000_0000 = 16384
        //
        // Products (float):
        // 0.5 * 2.0   = 1.0
        // 1.0 * 1.0   = 1.0
        // -0.5 * 1.0  = -0.5
        // 0.25 * 4.0  = 1.0
        // Sum = 2.5

        a0 = 16'b0010_0000_0000_0000; //  0.5
        b0 = 16'b0010_0000_0000_0000; //  2.0

        a1 = 16'b0100_0000_0000_0000; //  1.0
        b1 = 16'b0001_0000_0000_0000; //  1.0

        a2 = 16'b1110_0000_0000_0000; // -0.5
        b2 = 16'b0001_0000_0000_0000; //  1.0

        a3 = 16'b0001_0000_0000_0000; //  0.25
        b3 = 16'b0100_0000_0000_0000; //  4.0

        #1;

        // Expect 2.5 in Q4.12 = 2.5 * 4096 = 10240 = 0b_0010_1000_0000_0000
        if (result === 16'b0010_1000_0000_0000) begin
            $display("✅ PASS: result = %0d (Q4.12)", result);
        end else begin
            $display("❌ FAIL: result = %0d, expected 10240", result);
        end

        $finish;
    end

endmodule
